magic
tech sky130A
magscale 1 2
timestamp 1746697874
<< viali >>
rect 1593 8585 1627 8619
rect 3893 8585 3927 8619
rect 5365 8585 5399 8619
rect 7205 8585 7239 8619
rect 9045 8585 9079 8619
rect 10885 8585 10919 8619
rect 12725 8585 12759 8619
rect 14565 8585 14599 8619
rect 16773 8585 16807 8619
rect 18245 8585 18279 8619
rect 20085 8585 20119 8619
rect 21925 8585 21959 8619
rect 23765 8585 23799 8619
rect 25605 8585 25639 8619
rect 27445 8585 27479 8619
rect 29653 8585 29687 8619
rect 31125 8585 31159 8619
rect 32965 8585 32999 8619
rect 34805 8585 34839 8619
rect 36369 8585 36403 8619
rect 36645 8585 36679 8619
rect 38025 8585 38059 8619
rect 38393 8585 38427 8619
rect 1777 8449 1811 8483
rect 4077 8449 4111 8483
rect 5549 8449 5583 8483
rect 7389 8449 7423 8483
rect 9229 8449 9263 8483
rect 11069 8449 11103 8483
rect 12909 8449 12943 8483
rect 14749 8449 14783 8483
rect 16957 8449 16991 8483
rect 18429 8449 18463 8483
rect 20269 8449 20303 8483
rect 22109 8449 22143 8483
rect 23949 8449 23983 8483
rect 25789 8449 25823 8483
rect 27629 8449 27663 8483
rect 29837 8449 29871 8483
rect 31309 8449 31343 8483
rect 33149 8449 33183 8483
rect 34989 8449 35023 8483
rect 36185 8449 36219 8483
rect 36829 8449 36863 8483
rect 37473 8449 37507 8483
rect 37841 8449 37875 8483
rect 38209 8449 38243 8483
rect 37657 8313 37691 8347
rect 36921 8041 36955 8075
rect 37289 8041 37323 8075
rect 37657 8041 37691 8075
rect 36737 7837 36771 7871
rect 37105 7837 37139 7871
rect 37473 7837 37507 7871
rect 37841 7837 37875 7871
rect 38209 7837 38243 7871
rect 38025 7701 38059 7735
rect 38393 7701 38427 7735
rect 16405 7497 16439 7531
rect 16865 7497 16899 7531
rect 17049 7497 17083 7531
rect 17417 7497 17451 7531
rect 17693 7497 17727 7531
rect 18061 7497 18095 7531
rect 21833 7497 21867 7531
rect 22385 7497 22419 7531
rect 38025 7497 38059 7531
rect 16037 7429 16071 7463
rect 16497 7429 16531 7463
rect 15301 7361 15335 7395
rect 15485 7361 15519 7395
rect 15761 7361 15795 7395
rect 16313 7361 16347 7395
rect 16681 7361 16715 7395
rect 17233 7361 17267 7395
rect 17509 7361 17543 7395
rect 17969 7361 18003 7395
rect 18245 7361 18279 7395
rect 18613 7361 18647 7395
rect 19165 7361 19199 7395
rect 19257 7361 19291 7395
rect 19533 7361 19567 7395
rect 19809 7361 19843 7395
rect 20269 7361 20303 7395
rect 20545 7361 20579 7395
rect 20729 7361 20763 7395
rect 21557 7361 21591 7395
rect 22017 7361 22051 7395
rect 22569 7361 22603 7395
rect 23857 7361 23891 7395
rect 25421 7361 25455 7395
rect 25789 7361 25823 7395
rect 26249 7361 26283 7395
rect 26525 7361 26559 7395
rect 37841 7361 37875 7395
rect 38209 7361 38243 7395
rect 16221 7293 16255 7327
rect 17141 7293 17175 7327
rect 20453 7293 20487 7327
rect 15669 7225 15703 7259
rect 17785 7225 17819 7259
rect 18429 7225 18463 7259
rect 18797 7225 18831 7259
rect 19717 7225 19751 7259
rect 20729 7225 20763 7259
rect 21281 7225 21315 7259
rect 15945 7157 15979 7191
rect 18981 7157 19015 7191
rect 19993 7157 20027 7191
rect 20177 7157 20211 7191
rect 21373 7157 21407 7191
rect 23673 7157 23707 7191
rect 25237 7157 25271 7191
rect 25605 7157 25639 7191
rect 26065 7157 26099 7191
rect 26341 7157 26375 7191
rect 38393 7157 38427 7191
rect 15761 6817 15795 6851
rect 7389 6749 7423 6783
rect 7665 6749 7699 6783
rect 8125 6749 8159 6783
rect 8401 6749 8435 6783
rect 8953 6749 8987 6783
rect 9321 6749 9355 6783
rect 9873 6749 9907 6783
rect 10333 6749 10367 6783
rect 15853 6749 15887 6783
rect 15945 6749 15979 6783
rect 19993 6749 20027 6783
rect 26525 6749 26559 6783
rect 37841 6749 37875 6783
rect 38209 6749 38243 6783
rect 7573 6613 7607 6647
rect 7849 6613 7883 6647
rect 8309 6613 8343 6647
rect 8585 6613 8619 6647
rect 9137 6613 9171 6647
rect 9505 6613 9539 6647
rect 10057 6613 10091 6647
rect 10517 6613 10551 6647
rect 16129 6613 16163 6647
rect 20177 6613 20211 6647
rect 26341 6613 26375 6647
rect 38025 6613 38059 6647
rect 38393 6613 38427 6647
rect 9781 6409 9815 6443
rect 11161 6409 11195 6443
rect 16681 6409 16715 6443
rect 17049 6409 17083 6443
rect 38393 6409 38427 6443
rect 9597 6273 9631 6307
rect 10425 6273 10459 6307
rect 10977 6273 11011 6307
rect 16773 6273 16807 6307
rect 16865 6273 16899 6307
rect 37841 6273 37875 6307
rect 38209 6273 38243 6307
rect 10609 6137 10643 6171
rect 38025 6069 38059 6103
rect 18705 5865 18739 5899
rect 19073 5865 19107 5899
rect 28181 5865 28215 5899
rect 34253 5865 34287 5899
rect 35541 5865 35575 5899
rect 36737 5865 36771 5899
rect 37197 5865 37231 5899
rect 12817 5797 12851 5831
rect 14289 5797 14323 5831
rect 38393 5797 38427 5831
rect 21465 5729 21499 5763
rect 6009 5661 6043 5695
rect 7297 5661 7331 5695
rect 12633 5661 12667 5695
rect 12909 5661 12943 5695
rect 13185 5661 13219 5695
rect 13553 5661 13587 5695
rect 14105 5661 14139 5695
rect 18797 5661 18831 5695
rect 18889 5661 18923 5695
rect 21557 5661 21591 5695
rect 21649 5661 21683 5695
rect 28365 5661 28399 5695
rect 34437 5661 34471 5695
rect 35725 5661 35759 5695
rect 36921 5661 36955 5695
rect 37013 5661 37047 5695
rect 37841 5661 37875 5695
rect 38209 5661 38243 5695
rect 6193 5525 6227 5559
rect 7481 5525 7515 5559
rect 13093 5525 13127 5559
rect 13369 5525 13403 5559
rect 13737 5525 13771 5559
rect 21833 5525 21867 5559
rect 38025 5525 38059 5559
rect 4353 5321 4387 5355
rect 17417 5321 17451 5355
rect 17785 5321 17819 5355
rect 20177 5321 20211 5355
rect 23673 5321 23707 5355
rect 32873 5321 32907 5355
rect 38393 5321 38427 5355
rect 4169 5185 4203 5219
rect 4445 5185 4479 5219
rect 4721 5185 4755 5219
rect 5549 5185 5583 5219
rect 13737 5185 13771 5219
rect 14013 5185 14047 5219
rect 14289 5185 14323 5219
rect 14565 5185 14599 5219
rect 17509 5185 17543 5219
rect 17601 5185 17635 5219
rect 19809 5185 19843 5219
rect 19993 5185 20027 5219
rect 22937 5185 22971 5219
rect 23029 5185 23063 5219
rect 23397 5185 23431 5219
rect 23489 5185 23523 5219
rect 33057 5185 33091 5219
rect 37841 5185 37875 5219
rect 38209 5185 38243 5219
rect 14473 5049 14507 5083
rect 4629 4981 4663 5015
rect 4905 4981 4939 5015
rect 5733 4981 5767 5015
rect 13921 4981 13955 5015
rect 14197 4981 14231 5015
rect 14749 4981 14783 5015
rect 22845 4981 22879 5015
rect 23213 4981 23247 5015
rect 23305 4981 23339 5015
rect 38025 4981 38059 5015
rect 4445 4777 4479 4811
rect 15485 4777 15519 4811
rect 19349 4777 19383 4811
rect 19625 4777 19659 4811
rect 29561 4777 29595 4811
rect 30757 4777 30791 4811
rect 21741 4709 21775 4743
rect 28273 4709 28307 4743
rect 38393 4709 38427 4743
rect 4261 4573 4295 4607
rect 15025 4573 15059 4607
rect 15301 4573 15335 4607
rect 19349 4573 19383 4607
rect 19441 4573 19475 4607
rect 21373 4573 21407 4607
rect 21557 4573 21591 4607
rect 23581 4573 23615 4607
rect 27721 4549 27755 4583
rect 27997 4573 28031 4607
rect 28273 4573 28307 4607
rect 29009 4573 29043 4607
rect 29745 4573 29779 4607
rect 30941 4573 30975 4607
rect 37841 4573 37875 4607
rect 38209 4573 38243 4607
rect 23489 4505 23523 4539
rect 15209 4437 15243 4471
rect 23765 4437 23799 4471
rect 27629 4437 27663 4471
rect 27905 4437 27939 4471
rect 28181 4437 28215 4471
rect 28825 4437 28859 4471
rect 38025 4437 38059 4471
rect 2881 4097 2915 4131
rect 15945 4097 15979 4131
rect 19165 4097 19199 4131
rect 19257 4097 19291 4131
rect 21833 4097 21867 4131
rect 22109 4097 22143 4131
rect 25605 4097 25639 4131
rect 25697 4097 25731 4131
rect 26433 4097 26467 4131
rect 26525 4097 26559 4131
rect 27077 4097 27111 4131
rect 27721 4097 27755 4131
rect 28273 4097 28307 4131
rect 28365 4097 28399 4131
rect 28825 4097 28859 4131
rect 29101 4097 29135 4131
rect 29193 4097 29227 4131
rect 29469 4097 29503 4131
rect 29745 4097 29779 4131
rect 29837 4097 29871 4131
rect 30205 4097 30239 4131
rect 30481 4097 30515 4131
rect 30757 4097 30791 4131
rect 30849 4097 30883 4131
rect 31217 4097 31251 4131
rect 37841 4097 37875 4131
rect 38209 4097 38243 4131
rect 19073 4029 19107 4063
rect 30113 4029 30147 4063
rect 16129 3961 16163 3995
rect 22017 3961 22051 3995
rect 28089 3961 28123 3995
rect 28733 3961 28767 3995
rect 29377 3961 29411 3995
rect 38393 3961 38427 3995
rect 3065 3893 3099 3927
rect 19441 3893 19475 3927
rect 25513 3893 25547 3927
rect 25881 3893 25915 3927
rect 26433 3893 26467 3927
rect 26709 3893 26743 3927
rect 27261 3893 27295 3927
rect 27905 3893 27939 3927
rect 28549 3893 28583 3927
rect 28917 3893 28951 3927
rect 29653 3893 29687 3927
rect 30021 3893 30055 3927
rect 30297 3893 30331 3927
rect 30573 3893 30607 3927
rect 30849 3893 30883 3927
rect 31033 3893 31067 3927
rect 38025 3893 38059 3927
rect 17049 3689 17083 3723
rect 24869 3689 24903 3723
rect 16589 3621 16623 3655
rect 17693 3621 17727 3655
rect 21833 3621 21867 3655
rect 23581 3621 23615 3655
rect 23857 3621 23891 3655
rect 38393 3621 38427 3655
rect 3801 3485 3835 3519
rect 16405 3485 16439 3519
rect 16865 3485 16899 3519
rect 17509 3485 17543 3519
rect 17785 3485 17819 3519
rect 21005 3485 21039 3519
rect 21097 3485 21131 3519
rect 21649 3485 21683 3519
rect 22109 3485 22143 3519
rect 22569 3485 22603 3519
rect 22661 3485 22695 3519
rect 23121 3485 23155 3519
rect 23397 3485 23431 3519
rect 23673 3485 23707 3519
rect 23949 3485 23983 3519
rect 24409 3485 24443 3519
rect 24685 3485 24719 3519
rect 28825 3485 28859 3519
rect 29101 3485 29135 3519
rect 29285 3485 29319 3519
rect 29745 3485 29779 3519
rect 30021 3485 30055 3519
rect 30113 3485 30147 3519
rect 37841 3485 37875 3519
rect 38209 3485 38243 3519
rect 22477 3417 22511 3451
rect 23305 3417 23339 3451
rect 3985 3349 4019 3383
rect 17969 3349 18003 3383
rect 20913 3349 20947 3383
rect 21281 3349 21315 3383
rect 22293 3349 22327 3383
rect 22845 3349 22879 3383
rect 23029 3349 23063 3383
rect 23213 3349 23247 3383
rect 24133 3349 24167 3383
rect 24593 3349 24627 3383
rect 28733 3349 28767 3383
rect 28917 3349 28951 3383
rect 29561 3349 29595 3383
rect 29837 3349 29871 3383
rect 30205 3349 30239 3383
rect 38025 3349 38059 3383
rect 22569 3145 22603 3179
rect 38393 3145 38427 3179
rect 17509 3009 17543 3043
rect 18613 3009 18647 3043
rect 19441 3009 19475 3043
rect 22385 3009 22419 3043
rect 22753 3009 22787 3043
rect 23305 3009 23339 3043
rect 23857 3009 23891 3043
rect 24961 3009 24995 3043
rect 25789 3009 25823 3043
rect 26157 3009 26191 3043
rect 27445 3009 27479 3043
rect 28549 3009 28583 3043
rect 28917 3009 28951 3043
rect 29653 3009 29687 3043
rect 30481 3009 30515 3043
rect 31033 3009 31067 3043
rect 37473 3009 37507 3043
rect 37841 3009 37875 3043
rect 38209 3009 38243 3043
rect 26341 2873 26375 2907
rect 17693 2805 17727 2839
rect 18797 2805 18831 2839
rect 19625 2805 19659 2839
rect 22937 2805 22971 2839
rect 23489 2805 23523 2839
rect 24041 2805 24075 2839
rect 25145 2805 25179 2839
rect 25973 2805 26007 2839
rect 27261 2805 27295 2839
rect 28365 2805 28399 2839
rect 28733 2805 28767 2839
rect 29469 2805 29503 2839
rect 30665 2805 30699 2839
rect 31217 2805 31251 2839
rect 37657 2805 37691 2839
rect 38025 2805 38059 2839
rect 24593 2601 24627 2635
rect 25697 2601 25731 2635
rect 27905 2601 27939 2635
rect 28917 2601 28951 2635
rect 30849 2601 30883 2635
rect 22385 2533 22419 2567
rect 23121 2533 23155 2567
rect 24961 2533 24995 2567
rect 26065 2533 26099 2567
rect 27169 2533 27203 2567
rect 28273 2533 28307 2567
rect 29653 2533 29687 2567
rect 30481 2533 30515 2567
rect 31585 2533 31619 2567
rect 38393 2533 38427 2567
rect 16957 2397 16991 2431
rect 17325 2397 17359 2431
rect 17693 2397 17727 2431
rect 18061 2397 18095 2431
rect 18429 2397 18463 2431
rect 18797 2397 18831 2431
rect 19257 2397 19291 2431
rect 19625 2397 19659 2431
rect 19993 2397 20027 2431
rect 20361 2397 20395 2431
rect 20729 2397 20763 2431
rect 21097 2397 21131 2431
rect 21833 2397 21867 2431
rect 22201 2397 22235 2431
rect 22569 2397 22603 2431
rect 22937 2397 22971 2431
rect 23305 2397 23339 2431
rect 23673 2397 23707 2431
rect 24409 2397 24443 2431
rect 24777 2397 24811 2431
rect 25145 2397 25179 2431
rect 25513 2397 25547 2431
rect 25881 2397 25915 2431
rect 26249 2397 26283 2431
rect 26985 2397 27019 2431
rect 27353 2397 27387 2431
rect 27721 2397 27755 2431
rect 28089 2397 28123 2431
rect 28733 2397 28767 2431
rect 29101 2397 29135 2431
rect 29837 2397 29871 2431
rect 30205 2397 30239 2431
rect 30297 2397 30331 2431
rect 30665 2397 30699 2431
rect 31033 2397 31067 2431
rect 31401 2397 31435 2431
rect 32137 2397 32171 2431
rect 36461 2397 36495 2431
rect 36829 2397 36863 2431
rect 37473 2397 37507 2431
rect 37841 2397 37875 2431
rect 38209 2397 38243 2431
rect 17141 2261 17175 2295
rect 17509 2261 17543 2295
rect 17877 2261 17911 2295
rect 18245 2261 18279 2295
rect 18613 2261 18647 2295
rect 18981 2261 19015 2295
rect 19441 2261 19475 2295
rect 19809 2261 19843 2295
rect 20177 2261 20211 2295
rect 20545 2261 20579 2295
rect 20913 2261 20947 2295
rect 21281 2261 21315 2295
rect 22017 2261 22051 2295
rect 22753 2261 22787 2295
rect 23489 2261 23523 2295
rect 23857 2261 23891 2295
rect 25329 2261 25363 2295
rect 26433 2261 26467 2295
rect 27537 2261 27571 2295
rect 28549 2261 28583 2295
rect 30021 2261 30055 2295
rect 31217 2261 31251 2295
rect 32321 2261 32355 2295
rect 36645 2261 36679 2295
rect 37013 2261 37047 2295
rect 37657 2261 37691 2295
rect 38025 2261 38059 2295
<< metal1 >>
rect 7374 9256 7380 9308
rect 7432 9296 7438 9308
rect 20898 9296 20904 9308
rect 7432 9268 20904 9296
rect 7432 9256 7438 9268
rect 20898 9256 20904 9268
rect 20956 9256 20962 9308
rect 20346 9188 20352 9240
rect 20404 9228 20410 9240
rect 36170 9228 36176 9240
rect 20404 9200 36176 9228
rect 20404 9188 20410 9200
rect 36170 9188 36176 9200
rect 36228 9188 36234 9240
rect 14734 9120 14740 9172
rect 14792 9160 14798 9172
rect 23382 9160 23388 9172
rect 14792 9132 23388 9160
rect 14792 9120 14798 9132
rect 23382 9120 23388 9132
rect 23440 9120 23446 9172
rect 12894 9052 12900 9104
rect 12952 9092 12958 9104
rect 25130 9092 25136 9104
rect 12952 9064 25136 9092
rect 12952 9052 12958 9064
rect 25130 9052 25136 9064
rect 25188 9052 25194 9104
rect 17218 8984 17224 9036
rect 17276 9024 17282 9036
rect 23658 9024 23664 9036
rect 17276 8996 23664 9024
rect 17276 8984 17282 8996
rect 23658 8984 23664 8996
rect 23716 8984 23722 9036
rect 18506 8916 18512 8968
rect 18564 8956 18570 8968
rect 37826 8956 37832 8968
rect 18564 8928 37832 8956
rect 18564 8916 18570 8928
rect 37826 8916 37832 8928
rect 37884 8916 37890 8968
rect 5534 8848 5540 8900
rect 5592 8888 5598 8900
rect 16758 8888 16764 8900
rect 5592 8860 16764 8888
rect 5592 8848 5598 8860
rect 16758 8848 16764 8860
rect 16816 8848 16822 8900
rect 16942 8848 16948 8900
rect 17000 8888 17006 8900
rect 25866 8888 25872 8900
rect 17000 8860 25872 8888
rect 17000 8848 17006 8860
rect 25866 8848 25872 8860
rect 25924 8848 25930 8900
rect 10778 8780 10784 8832
rect 10836 8820 10842 8832
rect 16482 8820 16488 8832
rect 10836 8792 16488 8820
rect 10836 8780 10842 8792
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 18414 8780 18420 8832
rect 18472 8820 18478 8832
rect 26510 8820 26516 8832
rect 18472 8792 26516 8820
rect 18472 8780 18478 8792
rect 26510 8780 26516 8792
rect 26568 8780 26574 8832
rect 1104 8730 38824 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 9010 8730
rect 9062 8678 9074 8730
rect 9126 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 15010 8730
rect 15062 8678 15074 8730
rect 15126 8678 15138 8730
rect 15190 8678 15202 8730
rect 15254 8678 15266 8730
rect 15318 8678 21010 8730
rect 21062 8678 21074 8730
rect 21126 8678 21138 8730
rect 21190 8678 21202 8730
rect 21254 8678 21266 8730
rect 21318 8678 27010 8730
rect 27062 8678 27074 8730
rect 27126 8678 27138 8730
rect 27190 8678 27202 8730
rect 27254 8678 27266 8730
rect 27318 8678 33010 8730
rect 33062 8678 33074 8730
rect 33126 8678 33138 8730
rect 33190 8678 33202 8730
rect 33254 8678 33266 8730
rect 33318 8678 38824 8730
rect 1104 8656 38824 8678
rect 1486 8576 1492 8628
rect 1544 8616 1550 8628
rect 1581 8619 1639 8625
rect 1581 8616 1593 8619
rect 1544 8588 1593 8616
rect 1544 8576 1550 8588
rect 1581 8585 1593 8588
rect 1627 8585 1639 8619
rect 1581 8579 1639 8585
rect 3418 8576 3424 8628
rect 3476 8616 3482 8628
rect 3881 8619 3939 8625
rect 3881 8616 3893 8619
rect 3476 8588 3893 8616
rect 3476 8576 3482 8588
rect 3881 8585 3893 8588
rect 3927 8585 3939 8619
rect 3881 8579 3939 8585
rect 5166 8576 5172 8628
rect 5224 8616 5230 8628
rect 5353 8619 5411 8625
rect 5353 8616 5365 8619
rect 5224 8588 5365 8616
rect 5224 8576 5230 8588
rect 5353 8585 5365 8588
rect 5399 8585 5411 8619
rect 5353 8579 5411 8585
rect 7006 8576 7012 8628
rect 7064 8616 7070 8628
rect 7193 8619 7251 8625
rect 7193 8616 7205 8619
rect 7064 8588 7205 8616
rect 7064 8576 7070 8588
rect 7193 8585 7205 8588
rect 7239 8585 7251 8619
rect 7193 8579 7251 8585
rect 8846 8576 8852 8628
rect 8904 8616 8910 8628
rect 9033 8619 9091 8625
rect 9033 8616 9045 8619
rect 8904 8588 9045 8616
rect 8904 8576 8910 8588
rect 9033 8585 9045 8588
rect 9079 8585 9091 8619
rect 9033 8579 9091 8585
rect 10686 8576 10692 8628
rect 10744 8616 10750 8628
rect 10873 8619 10931 8625
rect 10873 8616 10885 8619
rect 10744 8588 10885 8616
rect 10744 8576 10750 8588
rect 10873 8585 10885 8588
rect 10919 8585 10931 8619
rect 10873 8579 10931 8585
rect 12526 8576 12532 8628
rect 12584 8616 12590 8628
rect 12713 8619 12771 8625
rect 12713 8616 12725 8619
rect 12584 8588 12725 8616
rect 12584 8576 12590 8588
rect 12713 8585 12725 8588
rect 12759 8585 12771 8619
rect 12713 8579 12771 8585
rect 14366 8576 14372 8628
rect 14424 8616 14430 8628
rect 14553 8619 14611 8625
rect 14553 8616 14565 8619
rect 14424 8588 14565 8616
rect 14424 8576 14430 8588
rect 14553 8585 14565 8588
rect 14599 8585 14611 8619
rect 14553 8579 14611 8585
rect 16206 8576 16212 8628
rect 16264 8616 16270 8628
rect 16761 8619 16819 8625
rect 16761 8616 16773 8619
rect 16264 8588 16773 8616
rect 16264 8576 16270 8588
rect 16761 8585 16773 8588
rect 16807 8585 16819 8619
rect 16761 8579 16819 8585
rect 18046 8576 18052 8628
rect 18104 8616 18110 8628
rect 18233 8619 18291 8625
rect 18233 8616 18245 8619
rect 18104 8588 18245 8616
rect 18104 8576 18110 8588
rect 18233 8585 18245 8588
rect 18279 8585 18291 8619
rect 18233 8579 18291 8585
rect 19886 8576 19892 8628
rect 19944 8616 19950 8628
rect 20073 8619 20131 8625
rect 20073 8616 20085 8619
rect 19944 8588 20085 8616
rect 19944 8576 19950 8588
rect 20073 8585 20085 8588
rect 20119 8585 20131 8619
rect 21634 8616 21640 8628
rect 20073 8579 20131 8585
rect 20180 8588 21640 8616
rect 17218 8548 17224 8560
rect 1780 8520 4292 8548
rect 1780 8489 1808 8520
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8449 1823 8483
rect 1765 8443 1823 8449
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 4080 8344 4108 8443
rect 4264 8412 4292 8520
rect 12406 8520 17224 8548
rect 5534 8440 5540 8492
rect 5592 8440 5598 8492
rect 7374 8440 7380 8492
rect 7432 8440 7438 8492
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8480 9275 8483
rect 10778 8480 10784 8492
rect 9263 8452 10784 8480
rect 9263 8449 9275 8452
rect 9217 8443 9275 8449
rect 10778 8440 10784 8452
rect 10836 8440 10842 8492
rect 11057 8483 11115 8489
rect 11057 8449 11069 8483
rect 11103 8480 11115 8483
rect 12406 8480 12434 8520
rect 17218 8508 17224 8520
rect 17276 8508 17282 8560
rect 17310 8508 17316 8560
rect 17368 8548 17374 8560
rect 20180 8548 20208 8588
rect 21634 8576 21640 8588
rect 21692 8576 21698 8628
rect 21726 8576 21732 8628
rect 21784 8616 21790 8628
rect 21913 8619 21971 8625
rect 21913 8616 21925 8619
rect 21784 8588 21925 8616
rect 21784 8576 21790 8588
rect 21913 8585 21925 8588
rect 21959 8585 21971 8619
rect 21913 8579 21971 8585
rect 23566 8576 23572 8628
rect 23624 8616 23630 8628
rect 23753 8619 23811 8625
rect 23753 8616 23765 8619
rect 23624 8588 23765 8616
rect 23624 8576 23630 8588
rect 23753 8585 23765 8588
rect 23799 8585 23811 8619
rect 23753 8579 23811 8585
rect 25406 8576 25412 8628
rect 25464 8616 25470 8628
rect 25593 8619 25651 8625
rect 25593 8616 25605 8619
rect 25464 8588 25605 8616
rect 25464 8576 25470 8588
rect 25593 8585 25605 8588
rect 25639 8585 25651 8619
rect 25593 8579 25651 8585
rect 27338 8576 27344 8628
rect 27396 8616 27402 8628
rect 27433 8619 27491 8625
rect 27433 8616 27445 8619
rect 27396 8588 27445 8616
rect 27396 8576 27402 8588
rect 27433 8585 27445 8588
rect 27479 8585 27491 8619
rect 27433 8579 27491 8585
rect 29086 8576 29092 8628
rect 29144 8616 29150 8628
rect 29641 8619 29699 8625
rect 29641 8616 29653 8619
rect 29144 8588 29653 8616
rect 29144 8576 29150 8588
rect 29641 8585 29653 8588
rect 29687 8585 29699 8619
rect 29641 8579 29699 8585
rect 30926 8576 30932 8628
rect 30984 8616 30990 8628
rect 31113 8619 31171 8625
rect 31113 8616 31125 8619
rect 30984 8588 31125 8616
rect 30984 8576 30990 8588
rect 31113 8585 31125 8588
rect 31159 8585 31171 8619
rect 31113 8579 31171 8585
rect 32766 8576 32772 8628
rect 32824 8616 32830 8628
rect 32953 8619 33011 8625
rect 32953 8616 32965 8619
rect 32824 8588 32965 8616
rect 32824 8576 32830 8588
rect 32953 8585 32965 8588
rect 32999 8585 33011 8619
rect 32953 8579 33011 8585
rect 34606 8576 34612 8628
rect 34664 8616 34670 8628
rect 34793 8619 34851 8625
rect 34793 8616 34805 8619
rect 34664 8588 34805 8616
rect 34664 8576 34670 8588
rect 34793 8585 34805 8588
rect 34839 8585 34851 8619
rect 34793 8579 34851 8585
rect 36354 8576 36360 8628
rect 36412 8576 36418 8628
rect 36446 8576 36452 8628
rect 36504 8616 36510 8628
rect 36633 8619 36691 8625
rect 36633 8616 36645 8619
rect 36504 8588 36645 8616
rect 36504 8576 36510 8588
rect 36633 8585 36645 8588
rect 36679 8585 36691 8619
rect 36633 8579 36691 8585
rect 38013 8619 38071 8625
rect 38013 8585 38025 8619
rect 38059 8585 38071 8619
rect 38013 8579 38071 8585
rect 25682 8548 25688 8560
rect 17368 8520 20208 8548
rect 20272 8520 25688 8548
rect 17368 8508 17374 8520
rect 11103 8452 12434 8480
rect 11103 8449 11115 8452
rect 11057 8443 11115 8449
rect 12894 8440 12900 8492
rect 12952 8440 12958 8492
rect 14734 8440 14740 8492
rect 14792 8440 14798 8492
rect 16942 8440 16948 8492
rect 17000 8440 17006 8492
rect 18414 8440 18420 8492
rect 18472 8440 18478 8492
rect 20272 8489 20300 8520
rect 25682 8508 25688 8520
rect 25740 8508 25746 8560
rect 38028 8548 38056 8579
rect 38286 8576 38292 8628
rect 38344 8616 38350 8628
rect 38381 8619 38439 8625
rect 38381 8616 38393 8619
rect 38344 8588 38393 8616
rect 38344 8576 38350 8588
rect 38381 8585 38393 8588
rect 38427 8585 38439 8619
rect 38381 8579 38439 8585
rect 38930 8548 38936 8560
rect 38028 8520 38936 8548
rect 38930 8508 38936 8520
rect 38988 8508 38994 8560
rect 20257 8483 20315 8489
rect 18524 8452 19656 8480
rect 18524 8412 18552 8452
rect 4264 8384 18552 8412
rect 19628 8412 19656 8452
rect 20257 8449 20269 8483
rect 20303 8449 20315 8483
rect 20257 8443 20315 8449
rect 22094 8440 22100 8492
rect 22152 8440 22158 8492
rect 23937 8483 23995 8489
rect 23937 8449 23949 8483
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 22370 8412 22376 8424
rect 19628 8384 22376 8412
rect 22370 8372 22376 8384
rect 22428 8372 22434 8424
rect 23952 8412 23980 8443
rect 25774 8440 25780 8492
rect 25832 8440 25838 8492
rect 27614 8440 27620 8492
rect 27672 8440 27678 8492
rect 29825 8483 29883 8489
rect 29825 8449 29837 8483
rect 29871 8480 29883 8483
rect 30742 8480 30748 8492
rect 29871 8452 30748 8480
rect 29871 8449 29883 8452
rect 29825 8443 29883 8449
rect 30742 8440 30748 8452
rect 30800 8440 30806 8492
rect 31294 8440 31300 8492
rect 31352 8440 31358 8492
rect 33137 8483 33195 8489
rect 33137 8449 33149 8483
rect 33183 8480 33195 8483
rect 34238 8480 34244 8492
rect 33183 8452 34244 8480
rect 33183 8449 33195 8452
rect 33137 8443 33195 8449
rect 34238 8440 34244 8452
rect 34296 8440 34302 8492
rect 34974 8440 34980 8492
rect 35032 8440 35038 8492
rect 36170 8440 36176 8492
rect 36228 8440 36234 8492
rect 36814 8440 36820 8492
rect 36872 8440 36878 8492
rect 37461 8483 37519 8489
rect 37461 8449 37473 8483
rect 37507 8449 37519 8483
rect 37461 8443 37519 8449
rect 28810 8412 28816 8424
rect 23952 8384 28816 8412
rect 28810 8372 28816 8384
rect 28868 8372 28874 8424
rect 17310 8344 17316 8356
rect 4080 8316 17316 8344
rect 17310 8304 17316 8316
rect 17368 8304 17374 8356
rect 19702 8304 19708 8356
rect 19760 8344 19766 8356
rect 37476 8344 37504 8443
rect 37826 8440 37832 8492
rect 37884 8440 37890 8492
rect 38197 8483 38255 8489
rect 38197 8449 38209 8483
rect 38243 8449 38255 8483
rect 38197 8443 38255 8449
rect 37550 8372 37556 8424
rect 37608 8412 37614 8424
rect 38212 8412 38240 8443
rect 37608 8384 38240 8412
rect 37608 8372 37614 8384
rect 19760 8316 37504 8344
rect 37645 8347 37703 8353
rect 19760 8304 19766 8316
rect 37645 8313 37657 8347
rect 37691 8344 37703 8347
rect 38746 8344 38752 8356
rect 37691 8316 38752 8344
rect 37691 8313 37703 8316
rect 37645 8307 37703 8313
rect 38746 8304 38752 8316
rect 38804 8304 38810 8356
rect 1104 8186 38824 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 13950 8186
rect 14002 8134 14014 8186
rect 14066 8134 14078 8186
rect 14130 8134 14142 8186
rect 14194 8134 14206 8186
rect 14258 8134 19950 8186
rect 20002 8134 20014 8186
rect 20066 8134 20078 8186
rect 20130 8134 20142 8186
rect 20194 8134 20206 8186
rect 20258 8134 25950 8186
rect 26002 8134 26014 8186
rect 26066 8134 26078 8186
rect 26130 8134 26142 8186
rect 26194 8134 26206 8186
rect 26258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 37950 8186
rect 38002 8134 38014 8186
rect 38066 8134 38078 8186
rect 38130 8134 38142 8186
rect 38194 8134 38206 8186
rect 38258 8134 38824 8186
rect 1104 8112 38824 8134
rect 36906 8032 36912 8084
rect 36964 8032 36970 8084
rect 37274 8032 37280 8084
rect 37332 8032 37338 8084
rect 37642 8032 37648 8084
rect 37700 8032 37706 8084
rect 25222 7964 25228 8016
rect 25280 8004 25286 8016
rect 26878 8004 26884 8016
rect 25280 7976 26884 8004
rect 25280 7964 25286 7976
rect 26878 7964 26884 7976
rect 26936 7964 26942 8016
rect 16850 7896 16856 7948
rect 16908 7936 16914 7948
rect 16908 7908 31754 7936
rect 16908 7896 16914 7908
rect 15654 7828 15660 7880
rect 15712 7868 15718 7880
rect 31726 7868 31754 7908
rect 36725 7871 36783 7877
rect 36725 7868 36737 7871
rect 15712 7840 25452 7868
rect 31726 7840 36737 7868
rect 15712 7828 15718 7840
rect 17678 7760 17684 7812
rect 17736 7800 17742 7812
rect 18690 7800 18696 7812
rect 17736 7772 18696 7800
rect 17736 7760 17742 7772
rect 18690 7760 18696 7772
rect 18748 7760 18754 7812
rect 18782 7760 18788 7812
rect 18840 7800 18846 7812
rect 25424 7800 25452 7840
rect 36725 7837 36737 7840
rect 36771 7837 36783 7871
rect 36725 7831 36783 7837
rect 37090 7828 37096 7880
rect 37148 7828 37154 7880
rect 37458 7828 37464 7880
rect 37516 7828 37522 7880
rect 37829 7871 37887 7877
rect 37829 7837 37841 7871
rect 37875 7837 37887 7871
rect 38197 7871 38255 7877
rect 38197 7868 38209 7871
rect 37829 7831 37887 7837
rect 37936 7840 38209 7868
rect 37844 7800 37872 7831
rect 18840 7772 25360 7800
rect 25424 7772 37872 7800
rect 18840 7760 18846 7772
rect 18230 7692 18236 7744
rect 18288 7732 18294 7744
rect 19242 7732 19248 7744
rect 18288 7704 19248 7732
rect 18288 7692 18294 7704
rect 19242 7692 19248 7704
rect 19300 7692 19306 7744
rect 20530 7692 20536 7744
rect 20588 7732 20594 7744
rect 25222 7732 25228 7744
rect 20588 7704 25228 7732
rect 20588 7692 20594 7704
rect 25222 7692 25228 7704
rect 25280 7692 25286 7744
rect 25332 7732 25360 7772
rect 37936 7732 37964 7840
rect 38197 7837 38209 7840
rect 38243 7837 38255 7871
rect 38197 7831 38255 7837
rect 25332 7704 37964 7732
rect 38010 7692 38016 7744
rect 38068 7692 38074 7744
rect 38378 7692 38384 7744
rect 38436 7692 38442 7744
rect 1104 7642 38824 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 9010 7642
rect 9062 7590 9074 7642
rect 9126 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 15010 7642
rect 15062 7590 15074 7642
rect 15126 7590 15138 7642
rect 15190 7590 15202 7642
rect 15254 7590 15266 7642
rect 15318 7590 21010 7642
rect 21062 7590 21074 7642
rect 21126 7590 21138 7642
rect 21190 7590 21202 7642
rect 21254 7590 21266 7642
rect 21318 7590 27010 7642
rect 27062 7590 27074 7642
rect 27126 7590 27138 7642
rect 27190 7590 27202 7642
rect 27254 7590 27266 7642
rect 27318 7590 33010 7642
rect 33062 7590 33074 7642
rect 33126 7590 33138 7642
rect 33190 7590 33202 7642
rect 33254 7590 33266 7642
rect 33318 7590 38824 7642
rect 1104 7568 38824 7590
rect 14918 7488 14924 7540
rect 14976 7528 14982 7540
rect 16393 7531 16451 7537
rect 16393 7528 16405 7531
rect 14976 7500 16405 7528
rect 14976 7488 14982 7500
rect 16393 7497 16405 7500
rect 16439 7497 16451 7531
rect 16393 7491 16451 7497
rect 16850 7488 16856 7540
rect 16908 7488 16914 7540
rect 17034 7488 17040 7540
rect 17092 7488 17098 7540
rect 17405 7531 17463 7537
rect 17405 7497 17417 7531
rect 17451 7497 17463 7531
rect 17405 7491 17463 7497
rect 14826 7420 14832 7472
rect 14884 7460 14890 7472
rect 16025 7463 16083 7469
rect 16025 7460 16037 7463
rect 14884 7432 16037 7460
rect 14884 7420 14890 7432
rect 15286 7352 15292 7404
rect 15344 7392 15350 7404
rect 15764 7401 15792 7432
rect 16025 7429 16037 7432
rect 16071 7429 16083 7463
rect 16025 7423 16083 7429
rect 16485 7463 16543 7469
rect 16485 7429 16497 7463
rect 16531 7460 16543 7463
rect 17420 7460 17448 7491
rect 17678 7488 17684 7540
rect 17736 7488 17742 7540
rect 18046 7488 18052 7540
rect 18104 7488 18110 7540
rect 18432 7500 21772 7528
rect 18432 7460 18460 7500
rect 16531 7432 17264 7460
rect 17420 7432 18460 7460
rect 16531 7429 16543 7432
rect 16485 7423 16543 7429
rect 17236 7401 17264 7432
rect 18690 7420 18696 7472
rect 18748 7460 18754 7472
rect 18748 7432 21680 7460
rect 18748 7420 18754 7432
rect 15473 7395 15531 7401
rect 15473 7392 15485 7395
rect 15344 7364 15485 7392
rect 15344 7352 15350 7364
rect 15473 7361 15485 7364
rect 15519 7361 15531 7395
rect 15473 7355 15531 7361
rect 15749 7395 15807 7401
rect 15749 7361 15761 7395
rect 15795 7361 15807 7395
rect 15749 7355 15807 7361
rect 16301 7395 16359 7401
rect 16301 7361 16313 7395
rect 16347 7392 16359 7395
rect 16669 7395 16727 7401
rect 16669 7392 16681 7395
rect 16347 7364 16681 7392
rect 16347 7361 16359 7364
rect 16301 7355 16359 7361
rect 16669 7361 16681 7364
rect 16715 7361 16727 7395
rect 16669 7355 16727 7361
rect 17221 7395 17279 7401
rect 17221 7361 17233 7395
rect 17267 7361 17279 7395
rect 17221 7355 17279 7361
rect 17497 7395 17555 7401
rect 17497 7361 17509 7395
rect 17543 7361 17555 7395
rect 17497 7355 17555 7361
rect 17957 7395 18015 7401
rect 17957 7361 17969 7395
rect 18003 7361 18015 7395
rect 17957 7355 18015 7361
rect 14642 7284 14648 7336
rect 14700 7324 14706 7336
rect 16209 7327 16267 7333
rect 16209 7324 16221 7327
rect 14700 7296 16221 7324
rect 14700 7284 14706 7296
rect 16209 7293 16221 7296
rect 16255 7293 16267 7327
rect 16209 7287 16267 7293
rect 17129 7327 17187 7333
rect 17129 7293 17141 7327
rect 17175 7324 17187 7327
rect 17512 7324 17540 7355
rect 17175 7296 17540 7324
rect 17175 7293 17187 7296
rect 17129 7287 17187 7293
rect 15654 7216 15660 7268
rect 15712 7216 15718 7268
rect 16482 7216 16488 7268
rect 16540 7256 16546 7268
rect 17773 7259 17831 7265
rect 17773 7256 17785 7259
rect 16540 7228 17785 7256
rect 16540 7216 16546 7228
rect 17773 7225 17785 7228
rect 17819 7225 17831 7259
rect 17972 7256 18000 7355
rect 18230 7352 18236 7404
rect 18288 7352 18294 7404
rect 18506 7392 18512 7404
rect 18432 7364 18512 7392
rect 18322 7256 18328 7268
rect 17972 7228 18328 7256
rect 17773 7219 17831 7225
rect 18322 7216 18328 7228
rect 18380 7216 18386 7268
rect 18432 7265 18460 7364
rect 18506 7352 18512 7364
rect 18564 7352 18570 7404
rect 18598 7352 18604 7404
rect 18656 7352 18662 7404
rect 19153 7395 19211 7401
rect 19153 7361 19165 7395
rect 19199 7361 19211 7395
rect 19153 7355 19211 7361
rect 19168 7324 19196 7355
rect 19242 7352 19248 7404
rect 19300 7352 19306 7404
rect 19518 7352 19524 7404
rect 19576 7352 19582 7404
rect 19794 7352 19800 7404
rect 19852 7392 19858 7404
rect 20257 7395 20315 7401
rect 20257 7392 20269 7395
rect 19852 7364 20269 7392
rect 19852 7352 19858 7364
rect 20257 7361 20269 7364
rect 20303 7361 20315 7395
rect 20257 7355 20315 7361
rect 20530 7352 20536 7404
rect 20588 7352 20594 7404
rect 20717 7395 20775 7401
rect 20717 7361 20729 7395
rect 20763 7392 20775 7395
rect 21358 7392 21364 7404
rect 20763 7364 21364 7392
rect 20763 7361 20775 7364
rect 20717 7355 20775 7361
rect 21358 7352 21364 7364
rect 21416 7352 21422 7404
rect 21545 7395 21603 7401
rect 21545 7392 21557 7395
rect 21468 7364 21557 7392
rect 20441 7327 20499 7333
rect 20441 7324 20453 7327
rect 18708 7296 18920 7324
rect 19168 7296 20453 7324
rect 18417 7259 18475 7265
rect 18417 7225 18429 7259
rect 18463 7225 18475 7259
rect 18417 7219 18475 7225
rect 18506 7216 18512 7268
rect 18564 7256 18570 7268
rect 18708 7256 18736 7296
rect 18564 7228 18736 7256
rect 18564 7216 18570 7228
rect 18782 7216 18788 7268
rect 18840 7216 18846 7268
rect 18892 7256 18920 7296
rect 20441 7293 20453 7296
rect 20487 7293 20499 7327
rect 20441 7287 20499 7293
rect 21468 7268 21496 7364
rect 21545 7361 21557 7364
rect 21591 7361 21603 7395
rect 21545 7355 21603 7361
rect 18892 7228 19656 7256
rect 15930 7148 15936 7200
rect 15988 7148 15994 7200
rect 16758 7148 16764 7200
rect 16816 7188 16822 7200
rect 18969 7191 19027 7197
rect 18969 7188 18981 7191
rect 16816 7160 18981 7188
rect 16816 7148 16822 7160
rect 18969 7157 18981 7160
rect 19015 7157 19027 7191
rect 19628 7188 19656 7228
rect 19702 7216 19708 7268
rect 19760 7216 19766 7268
rect 20717 7259 20775 7265
rect 20717 7256 20729 7259
rect 19904 7228 20729 7256
rect 19904 7188 19932 7228
rect 20717 7225 20729 7228
rect 20763 7225 20775 7259
rect 20717 7219 20775 7225
rect 21269 7259 21327 7265
rect 21269 7225 21281 7259
rect 21315 7256 21327 7259
rect 21450 7256 21456 7268
rect 21315 7228 21456 7256
rect 21315 7225 21327 7228
rect 21269 7219 21327 7225
rect 21450 7216 21456 7228
rect 21508 7216 21514 7268
rect 21652 7256 21680 7432
rect 21744 7324 21772 7500
rect 21818 7488 21824 7540
rect 21876 7488 21882 7540
rect 22370 7488 22376 7540
rect 22428 7488 22434 7540
rect 32582 7528 32588 7540
rect 23308 7500 32588 7528
rect 23308 7460 23336 7500
rect 32582 7488 32588 7500
rect 32640 7488 32646 7540
rect 38013 7531 38071 7537
rect 38013 7497 38025 7531
rect 38059 7528 38071 7531
rect 38470 7528 38476 7540
rect 38059 7500 38476 7528
rect 38059 7497 38071 7500
rect 38013 7491 38071 7497
rect 38470 7488 38476 7500
rect 38528 7488 38534 7540
rect 21836 7432 23336 7460
rect 21836 7404 21864 7432
rect 23382 7420 23388 7472
rect 23440 7460 23446 7472
rect 25314 7460 25320 7472
rect 23440 7432 25320 7460
rect 23440 7420 23446 7432
rect 25314 7420 25320 7432
rect 25372 7420 25378 7472
rect 26142 7460 26148 7472
rect 25424 7432 26148 7460
rect 21818 7352 21824 7404
rect 21876 7352 21882 7404
rect 22005 7395 22063 7401
rect 22005 7361 22017 7395
rect 22051 7392 22063 7395
rect 22278 7392 22284 7404
rect 22051 7364 22284 7392
rect 22051 7361 22063 7364
rect 22005 7355 22063 7361
rect 22278 7352 22284 7364
rect 22336 7352 22342 7404
rect 22554 7352 22560 7404
rect 22612 7352 22618 7404
rect 23845 7395 23903 7401
rect 23845 7361 23857 7395
rect 23891 7392 23903 7395
rect 24118 7392 24124 7404
rect 23891 7364 24124 7392
rect 23891 7361 23903 7364
rect 23845 7355 23903 7361
rect 24118 7352 24124 7364
rect 24176 7352 24182 7404
rect 25424 7401 25452 7432
rect 26142 7420 26148 7432
rect 26200 7420 26206 7472
rect 26418 7420 26424 7472
rect 26476 7460 26482 7472
rect 26476 7432 37872 7460
rect 26476 7420 26482 7432
rect 25409 7395 25467 7401
rect 25409 7361 25421 7395
rect 25455 7361 25467 7395
rect 25409 7355 25467 7361
rect 25590 7352 25596 7404
rect 25648 7392 25654 7404
rect 25777 7395 25835 7401
rect 25777 7392 25789 7395
rect 25648 7364 25789 7392
rect 25648 7352 25654 7364
rect 25777 7361 25789 7364
rect 25823 7361 25835 7395
rect 25777 7355 25835 7361
rect 26237 7395 26295 7401
rect 26237 7361 26249 7395
rect 26283 7361 26295 7395
rect 26237 7355 26295 7361
rect 26513 7395 26571 7401
rect 26513 7361 26525 7395
rect 26559 7392 26571 7395
rect 33962 7392 33968 7404
rect 26559 7364 33968 7392
rect 26559 7361 26571 7364
rect 26513 7355 26571 7361
rect 26142 7324 26148 7336
rect 21744 7296 26148 7324
rect 26142 7284 26148 7296
rect 26200 7284 26206 7336
rect 26252 7324 26280 7355
rect 33962 7352 33968 7364
rect 34020 7352 34026 7404
rect 37844 7401 37872 7432
rect 37829 7395 37887 7401
rect 37829 7361 37841 7395
rect 37875 7361 37887 7395
rect 37829 7355 37887 7361
rect 38197 7395 38255 7401
rect 38197 7361 38209 7395
rect 38243 7361 38255 7395
rect 38197 7355 38255 7361
rect 26602 7324 26608 7336
rect 26252 7296 26608 7324
rect 26602 7284 26608 7296
rect 26660 7284 26666 7336
rect 26878 7284 26884 7336
rect 26936 7324 26942 7336
rect 31846 7324 31852 7336
rect 26936 7296 31852 7324
rect 26936 7284 26942 7296
rect 31846 7284 31852 7296
rect 31904 7284 31910 7336
rect 37274 7284 37280 7336
rect 37332 7324 37338 7336
rect 38212 7324 38240 7355
rect 37332 7296 38240 7324
rect 37332 7284 37338 7296
rect 37458 7256 37464 7268
rect 21652 7228 37464 7256
rect 37458 7216 37464 7228
rect 37516 7216 37522 7268
rect 19628 7160 19932 7188
rect 19981 7191 20039 7197
rect 18969 7151 19027 7157
rect 19981 7157 19993 7191
rect 20027 7188 20039 7191
rect 20070 7188 20076 7200
rect 20027 7160 20076 7188
rect 20027 7157 20039 7160
rect 19981 7151 20039 7157
rect 20070 7148 20076 7160
rect 20128 7148 20134 7200
rect 20165 7191 20223 7197
rect 20165 7157 20177 7191
rect 20211 7188 20223 7191
rect 20254 7188 20260 7200
rect 20211 7160 20260 7188
rect 20211 7157 20223 7160
rect 20165 7151 20223 7157
rect 20254 7148 20260 7160
rect 20312 7148 20318 7200
rect 20898 7148 20904 7200
rect 20956 7188 20962 7200
rect 21361 7191 21419 7197
rect 21361 7188 21373 7191
rect 20956 7160 21373 7188
rect 20956 7148 20962 7160
rect 21361 7157 21373 7160
rect 21407 7157 21419 7191
rect 21361 7151 21419 7157
rect 23658 7148 23664 7200
rect 23716 7148 23722 7200
rect 25130 7148 25136 7200
rect 25188 7188 25194 7200
rect 25225 7191 25283 7197
rect 25225 7188 25237 7191
rect 25188 7160 25237 7188
rect 25188 7148 25194 7160
rect 25225 7157 25237 7160
rect 25271 7157 25283 7191
rect 25225 7151 25283 7157
rect 25314 7148 25320 7200
rect 25372 7188 25378 7200
rect 25593 7191 25651 7197
rect 25593 7188 25605 7191
rect 25372 7160 25605 7188
rect 25372 7148 25378 7160
rect 25593 7157 25605 7160
rect 25639 7157 25651 7191
rect 25593 7151 25651 7157
rect 25866 7148 25872 7200
rect 25924 7188 25930 7200
rect 26053 7191 26111 7197
rect 26053 7188 26065 7191
rect 25924 7160 26065 7188
rect 25924 7148 25930 7160
rect 26053 7157 26065 7160
rect 26099 7157 26111 7191
rect 26053 7151 26111 7157
rect 26329 7191 26387 7197
rect 26329 7157 26341 7191
rect 26375 7188 26387 7191
rect 26510 7188 26516 7200
rect 26375 7160 26516 7188
rect 26375 7157 26387 7160
rect 26329 7151 26387 7157
rect 26510 7148 26516 7160
rect 26568 7148 26574 7200
rect 38378 7148 38384 7200
rect 38436 7148 38442 7200
rect 1104 7098 38824 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 13950 7098
rect 14002 7046 14014 7098
rect 14066 7046 14078 7098
rect 14130 7046 14142 7098
rect 14194 7046 14206 7098
rect 14258 7046 19950 7098
rect 20002 7046 20014 7098
rect 20066 7046 20078 7098
rect 20130 7046 20142 7098
rect 20194 7046 20206 7098
rect 20258 7046 25950 7098
rect 26002 7046 26014 7098
rect 26066 7046 26078 7098
rect 26130 7046 26142 7098
rect 26194 7046 26206 7098
rect 26258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 37950 7098
rect 38002 7046 38014 7098
rect 38066 7046 38078 7098
rect 38130 7046 38142 7098
rect 38194 7046 38206 7098
rect 38258 7046 38824 7098
rect 1104 7024 38824 7046
rect 15930 6944 15936 6996
rect 15988 6984 15994 6996
rect 37090 6984 37096 6996
rect 15988 6956 37096 6984
rect 15988 6944 15994 6956
rect 37090 6944 37096 6956
rect 37148 6944 37154 6996
rect 7300 6888 7972 6916
rect 1302 6808 1308 6860
rect 1360 6848 1366 6860
rect 7300 6848 7328 6888
rect 7834 6848 7840 6860
rect 1360 6820 7328 6848
rect 7392 6820 7840 6848
rect 1360 6808 1366 6820
rect 7392 6789 7420 6820
rect 7834 6808 7840 6820
rect 7892 6808 7898 6860
rect 7944 6848 7972 6888
rect 7944 6820 12434 6848
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6749 7435 6783
rect 7377 6743 7435 6749
rect 7653 6783 7711 6789
rect 7653 6749 7665 6783
rect 7699 6780 7711 6783
rect 7742 6780 7748 6792
rect 7699 6752 7748 6780
rect 7699 6749 7711 6752
rect 7653 6743 7711 6749
rect 7742 6740 7748 6752
rect 7800 6740 7806 6792
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 7466 6672 7472 6724
rect 7524 6712 7530 6724
rect 8128 6712 8156 6743
rect 8386 6740 8392 6792
rect 8444 6740 8450 6792
rect 8941 6783 8999 6789
rect 8941 6749 8953 6783
rect 8987 6749 8999 6783
rect 9309 6783 9367 6789
rect 9309 6780 9321 6783
rect 8941 6743 8999 6749
rect 9048 6752 9321 6780
rect 7524 6684 8156 6712
rect 7524 6672 7530 6684
rect 8202 6672 8208 6724
rect 8260 6712 8266 6724
rect 8956 6712 8984 6743
rect 8260 6684 8984 6712
rect 8260 6672 8266 6684
rect 7558 6604 7564 6656
rect 7616 6604 7622 6656
rect 7650 6604 7656 6656
rect 7708 6644 7714 6656
rect 7837 6647 7895 6653
rect 7837 6644 7849 6647
rect 7708 6616 7849 6644
rect 7708 6604 7714 6616
rect 7837 6613 7849 6616
rect 7883 6613 7895 6647
rect 7837 6607 7895 6613
rect 8297 6647 8355 6653
rect 8297 6613 8309 6647
rect 8343 6644 8355 6647
rect 8478 6644 8484 6656
rect 8343 6616 8484 6644
rect 8343 6613 8355 6616
rect 8297 6607 8355 6613
rect 8478 6604 8484 6616
rect 8536 6604 8542 6656
rect 8570 6604 8576 6656
rect 8628 6604 8634 6656
rect 8662 6604 8668 6656
rect 8720 6644 8726 6656
rect 9048 6644 9076 6752
rect 9309 6749 9321 6752
rect 9355 6749 9367 6783
rect 9309 6743 9367 6749
rect 9490 6740 9496 6792
rect 9548 6780 9554 6792
rect 9861 6783 9919 6789
rect 9861 6780 9873 6783
rect 9548 6752 9873 6780
rect 9548 6740 9554 6752
rect 9861 6749 9873 6752
rect 9907 6749 9919 6783
rect 9861 6743 9919 6749
rect 10318 6740 10324 6792
rect 10376 6740 10382 6792
rect 11790 6712 11796 6724
rect 10060 6684 11796 6712
rect 8720 6616 9076 6644
rect 9125 6647 9183 6653
rect 8720 6604 8726 6616
rect 9125 6613 9137 6647
rect 9171 6644 9183 6647
rect 9398 6644 9404 6656
rect 9171 6616 9404 6644
rect 9171 6613 9183 6616
rect 9125 6607 9183 6613
rect 9398 6604 9404 6616
rect 9456 6604 9462 6656
rect 9493 6647 9551 6653
rect 9493 6613 9505 6647
rect 9539 6644 9551 6647
rect 9950 6644 9956 6656
rect 9539 6616 9956 6644
rect 9539 6613 9551 6616
rect 9493 6607 9551 6613
rect 9950 6604 9956 6616
rect 10008 6604 10014 6656
rect 10060 6653 10088 6684
rect 11790 6672 11796 6684
rect 11848 6672 11854 6724
rect 12406 6712 12434 6820
rect 15746 6808 15752 6860
rect 15804 6808 15810 6860
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6780 15899 6783
rect 15933 6783 15991 6789
rect 15933 6780 15945 6783
rect 15887 6752 15945 6780
rect 15887 6749 15899 6752
rect 15841 6743 15899 6749
rect 15933 6749 15945 6752
rect 15979 6749 15991 6783
rect 15933 6743 15991 6749
rect 19981 6783 20039 6789
rect 19981 6749 19993 6783
rect 20027 6749 20039 6783
rect 19981 6743 20039 6749
rect 26513 6783 26571 6789
rect 26513 6749 26525 6783
rect 26559 6780 26571 6783
rect 34146 6780 34152 6792
rect 26559 6752 34152 6780
rect 26559 6749 26571 6752
rect 26513 6743 26571 6749
rect 19996 6712 20024 6743
rect 34146 6740 34152 6752
rect 34204 6740 34210 6792
rect 37829 6783 37887 6789
rect 37829 6749 37841 6783
rect 37875 6749 37887 6783
rect 37829 6743 37887 6749
rect 12406 6684 20024 6712
rect 20070 6672 20076 6724
rect 20128 6712 20134 6724
rect 37844 6712 37872 6743
rect 38194 6740 38200 6792
rect 38252 6740 38258 6792
rect 20128 6684 37872 6712
rect 20128 6672 20134 6684
rect 10045 6647 10103 6653
rect 10045 6613 10057 6647
rect 10091 6613 10103 6647
rect 10045 6607 10103 6613
rect 10505 6647 10563 6653
rect 10505 6613 10517 6647
rect 10551 6644 10563 6647
rect 11606 6644 11612 6656
rect 10551 6616 11612 6644
rect 10551 6613 10563 6616
rect 10505 6607 10563 6613
rect 11606 6604 11612 6616
rect 11664 6604 11670 6656
rect 16114 6604 16120 6656
rect 16172 6604 16178 6656
rect 20162 6604 20168 6656
rect 20220 6604 20226 6656
rect 25682 6604 25688 6656
rect 25740 6644 25746 6656
rect 26329 6647 26387 6653
rect 26329 6644 26341 6647
rect 25740 6616 26341 6644
rect 25740 6604 25746 6616
rect 26329 6613 26341 6616
rect 26375 6613 26387 6647
rect 26329 6607 26387 6613
rect 38010 6604 38016 6656
rect 38068 6604 38074 6656
rect 38378 6604 38384 6656
rect 38436 6604 38442 6656
rect 1104 6554 38824 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 9010 6554
rect 9062 6502 9074 6554
rect 9126 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 15010 6554
rect 15062 6502 15074 6554
rect 15126 6502 15138 6554
rect 15190 6502 15202 6554
rect 15254 6502 15266 6554
rect 15318 6502 21010 6554
rect 21062 6502 21074 6554
rect 21126 6502 21138 6554
rect 21190 6502 21202 6554
rect 21254 6502 21266 6554
rect 21318 6502 27010 6554
rect 27062 6502 27074 6554
rect 27126 6502 27138 6554
rect 27190 6502 27202 6554
rect 27254 6502 27266 6554
rect 27318 6502 33010 6554
rect 33062 6502 33074 6554
rect 33126 6502 33138 6554
rect 33190 6502 33202 6554
rect 33254 6502 33266 6554
rect 33318 6502 38824 6554
rect 1104 6480 38824 6502
rect 6914 6400 6920 6452
rect 6972 6440 6978 6452
rect 8662 6440 8668 6452
rect 6972 6412 8668 6440
rect 6972 6400 6978 6412
rect 8662 6400 8668 6412
rect 8720 6400 8726 6452
rect 9769 6443 9827 6449
rect 9769 6409 9781 6443
rect 9815 6440 9827 6443
rect 10962 6440 10968 6452
rect 9815 6412 10968 6440
rect 9815 6409 9827 6412
rect 9769 6403 9827 6409
rect 10962 6400 10968 6412
rect 11020 6400 11026 6452
rect 11149 6443 11207 6449
rect 11149 6409 11161 6443
rect 11195 6409 11207 6443
rect 11149 6403 11207 6409
rect 7558 6332 7564 6384
rect 7616 6372 7622 6384
rect 11054 6372 11060 6384
rect 7616 6344 11060 6372
rect 7616 6332 7622 6344
rect 11054 6332 11060 6344
rect 11112 6332 11118 6384
rect 11164 6372 11192 6403
rect 16666 6400 16672 6452
rect 16724 6400 16730 6452
rect 17037 6443 17095 6449
rect 17037 6409 17049 6443
rect 17083 6440 17095 6443
rect 20070 6440 20076 6452
rect 17083 6412 20076 6440
rect 17083 6409 17095 6412
rect 17037 6403 17095 6409
rect 20070 6400 20076 6412
rect 20128 6400 20134 6452
rect 20162 6400 20168 6452
rect 20220 6440 20226 6452
rect 37274 6440 37280 6452
rect 20220 6412 37280 6440
rect 20220 6400 20226 6412
rect 37274 6400 37280 6412
rect 37332 6400 37338 6452
rect 38378 6400 38384 6452
rect 38436 6400 38442 6452
rect 15194 6372 15200 6384
rect 11164 6344 15200 6372
rect 15194 6332 15200 6344
rect 15252 6332 15258 6384
rect 19058 6332 19064 6384
rect 19116 6372 19122 6384
rect 19116 6344 38240 6372
rect 19116 6332 19122 6344
rect 6638 6264 6644 6316
rect 6696 6304 6702 6316
rect 9490 6304 9496 6316
rect 6696 6276 9496 6304
rect 6696 6264 6702 6276
rect 9490 6264 9496 6276
rect 9548 6264 9554 6316
rect 9582 6264 9588 6316
rect 9640 6264 9646 6316
rect 10413 6307 10471 6313
rect 10413 6273 10425 6307
rect 10459 6273 10471 6307
rect 10413 6267 10471 6273
rect 8294 6196 8300 6248
rect 8352 6236 8358 6248
rect 10428 6236 10456 6267
rect 10502 6264 10508 6316
rect 10560 6304 10566 6316
rect 10965 6307 11023 6313
rect 10965 6304 10977 6307
rect 10560 6276 10977 6304
rect 10560 6264 10566 6276
rect 10965 6273 10977 6276
rect 11011 6273 11023 6307
rect 10965 6267 11023 6273
rect 11330 6264 11336 6316
rect 11388 6304 11394 6316
rect 16574 6304 16580 6316
rect 11388 6276 16580 6304
rect 11388 6264 11394 6276
rect 16574 6264 16580 6276
rect 16632 6264 16638 6316
rect 16761 6307 16819 6313
rect 16761 6273 16773 6307
rect 16807 6304 16819 6307
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 16807 6276 16865 6304
rect 16807 6273 16819 6276
rect 16761 6267 16819 6273
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 17770 6264 17776 6316
rect 17828 6304 17834 6316
rect 38212 6313 38240 6344
rect 37829 6307 37887 6313
rect 37829 6304 37841 6307
rect 17828 6276 37841 6304
rect 17828 6264 17834 6276
rect 37829 6273 37841 6276
rect 37875 6273 37887 6307
rect 37829 6267 37887 6273
rect 38197 6307 38255 6313
rect 38197 6273 38209 6307
rect 38243 6273 38255 6307
rect 38197 6267 38255 6273
rect 8352 6208 10456 6236
rect 8352 6196 8358 6208
rect 11238 6196 11244 6248
rect 11296 6236 11302 6248
rect 18782 6236 18788 6248
rect 11296 6208 18788 6236
rect 11296 6196 11302 6208
rect 18782 6196 18788 6208
rect 18840 6196 18846 6248
rect 6086 6128 6092 6180
rect 6144 6168 6150 6180
rect 10502 6168 10508 6180
rect 6144 6140 10508 6168
rect 6144 6128 6150 6140
rect 10502 6128 10508 6140
rect 10560 6128 10566 6180
rect 10594 6128 10600 6180
rect 10652 6128 10658 6180
rect 11146 6128 11152 6180
rect 11204 6168 11210 6180
rect 18874 6168 18880 6180
rect 11204 6140 18880 6168
rect 11204 6128 11210 6140
rect 18874 6128 18880 6140
rect 18932 6128 18938 6180
rect 20346 6128 20352 6180
rect 20404 6168 20410 6180
rect 37826 6168 37832 6180
rect 20404 6140 37832 6168
rect 20404 6128 20410 6140
rect 37826 6128 37832 6140
rect 37884 6128 37890 6180
rect 7190 6060 7196 6112
rect 7248 6100 7254 6112
rect 8202 6100 8208 6112
rect 7248 6072 8208 6100
rect 7248 6060 7254 6072
rect 8202 6060 8208 6072
rect 8260 6060 8266 6112
rect 8570 6060 8576 6112
rect 8628 6100 8634 6112
rect 12618 6100 12624 6112
rect 8628 6072 12624 6100
rect 8628 6060 8634 6072
rect 12618 6060 12624 6072
rect 12676 6060 12682 6112
rect 12710 6060 12716 6112
rect 12768 6100 12774 6112
rect 19702 6100 19708 6112
rect 12768 6072 19708 6100
rect 12768 6060 12774 6072
rect 19702 6060 19708 6072
rect 19760 6060 19766 6112
rect 38013 6103 38071 6109
rect 38013 6069 38025 6103
rect 38059 6100 38071 6103
rect 39114 6100 39120 6112
rect 38059 6072 39120 6100
rect 38059 6069 38071 6072
rect 38013 6063 38071 6069
rect 39114 6060 39120 6072
rect 39172 6060 39178 6112
rect 1104 6010 38824 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 13950 6010
rect 14002 5958 14014 6010
rect 14066 5958 14078 6010
rect 14130 5958 14142 6010
rect 14194 5958 14206 6010
rect 14258 5958 19950 6010
rect 20002 5958 20014 6010
rect 20066 5958 20078 6010
rect 20130 5958 20142 6010
rect 20194 5958 20206 6010
rect 20258 5958 25950 6010
rect 26002 5958 26014 6010
rect 26066 5958 26078 6010
rect 26130 5958 26142 6010
rect 26194 5958 26206 6010
rect 26258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 37950 6010
rect 38002 5958 38014 6010
rect 38066 5958 38078 6010
rect 38130 5958 38142 6010
rect 38194 5958 38206 6010
rect 38258 5958 38824 6010
rect 1104 5936 38824 5958
rect 7650 5856 7656 5908
rect 7708 5896 7714 5908
rect 11146 5896 11152 5908
rect 7708 5868 11152 5896
rect 7708 5856 7714 5868
rect 11146 5856 11152 5868
rect 11204 5856 11210 5908
rect 18506 5896 18512 5908
rect 12544 5868 18512 5896
rect 6362 5788 6368 5840
rect 6420 5828 6426 5840
rect 10318 5828 10324 5840
rect 6420 5800 10324 5828
rect 6420 5788 6426 5800
rect 10318 5788 10324 5800
rect 10376 5788 10382 5840
rect 10594 5788 10600 5840
rect 10652 5828 10658 5840
rect 12544 5828 12572 5868
rect 18506 5856 18512 5868
rect 18564 5856 18570 5908
rect 18690 5856 18696 5908
rect 18748 5856 18754 5908
rect 19058 5856 19064 5908
rect 19116 5856 19122 5908
rect 22094 5856 22100 5908
rect 22152 5896 22158 5908
rect 28169 5899 28227 5905
rect 28169 5896 28181 5899
rect 22152 5868 28181 5896
rect 22152 5856 22158 5868
rect 28169 5865 28181 5868
rect 28215 5865 28227 5899
rect 28169 5859 28227 5865
rect 34238 5856 34244 5908
rect 34296 5856 34302 5908
rect 34974 5856 34980 5908
rect 35032 5896 35038 5908
rect 35529 5899 35587 5905
rect 35529 5896 35541 5899
rect 35032 5868 35541 5896
rect 35032 5856 35038 5868
rect 35529 5865 35541 5868
rect 35575 5865 35587 5899
rect 35529 5859 35587 5865
rect 36725 5899 36783 5905
rect 36725 5865 36737 5899
rect 36771 5896 36783 5899
rect 36814 5896 36820 5908
rect 36771 5868 36820 5896
rect 36771 5865 36783 5868
rect 36725 5859 36783 5865
rect 36814 5856 36820 5868
rect 36872 5856 36878 5908
rect 37185 5899 37243 5905
rect 37185 5865 37197 5899
rect 37231 5896 37243 5899
rect 37550 5896 37556 5908
rect 37231 5868 37556 5896
rect 37231 5865 37243 5868
rect 37185 5859 37243 5865
rect 37550 5856 37556 5868
rect 37608 5856 37614 5908
rect 10652 5800 12572 5828
rect 12805 5831 12863 5837
rect 10652 5788 10658 5800
rect 12805 5797 12817 5831
rect 12851 5828 12863 5831
rect 12851 5800 14228 5828
rect 12851 5797 12863 5800
rect 12805 5791 12863 5797
rect 4154 5720 4160 5772
rect 4212 5760 4218 5772
rect 9582 5760 9588 5772
rect 4212 5732 9588 5760
rect 4212 5720 4218 5732
rect 9582 5720 9588 5732
rect 9640 5720 9646 5772
rect 11054 5720 11060 5772
rect 11112 5760 11118 5772
rect 14200 5760 14228 5800
rect 14274 5788 14280 5840
rect 14332 5788 14338 5840
rect 15194 5788 15200 5840
rect 15252 5828 15258 5840
rect 22922 5828 22928 5840
rect 15252 5800 22928 5828
rect 15252 5788 15258 5800
rect 22922 5788 22928 5800
rect 22980 5788 22986 5840
rect 34514 5828 34520 5840
rect 31726 5800 34520 5828
rect 19334 5760 19340 5772
rect 11112 5732 12940 5760
rect 14200 5732 19340 5760
rect 11112 5720 11118 5732
rect 4982 5652 4988 5704
rect 5040 5692 5046 5704
rect 5997 5695 6055 5701
rect 5997 5692 6009 5695
rect 5040 5664 6009 5692
rect 5040 5652 5046 5664
rect 5997 5661 6009 5664
rect 6043 5661 6055 5695
rect 5997 5655 6055 5661
rect 7285 5695 7343 5701
rect 7285 5661 7297 5695
rect 7331 5661 7343 5695
rect 7285 5655 7343 5661
rect 4706 5584 4712 5636
rect 4764 5624 4770 5636
rect 7300 5624 7328 5655
rect 11422 5652 11428 5704
rect 11480 5692 11486 5704
rect 12912 5701 12940 5732
rect 19334 5720 19340 5732
rect 19392 5720 19398 5772
rect 21358 5720 21364 5772
rect 21416 5760 21422 5772
rect 21453 5763 21511 5769
rect 21453 5760 21465 5763
rect 21416 5732 21465 5760
rect 21416 5720 21422 5732
rect 21453 5729 21465 5732
rect 21499 5729 21511 5763
rect 21453 5723 21511 5729
rect 12621 5695 12679 5701
rect 12621 5692 12633 5695
rect 11480 5664 12633 5692
rect 11480 5652 11486 5664
rect 12621 5661 12633 5664
rect 12667 5661 12679 5695
rect 12621 5655 12679 5661
rect 12897 5695 12955 5701
rect 12897 5661 12909 5695
rect 12943 5661 12955 5695
rect 12897 5655 12955 5661
rect 13170 5652 13176 5704
rect 13228 5652 13234 5704
rect 13538 5652 13544 5704
rect 13596 5652 13602 5704
rect 13630 5652 13636 5704
rect 13688 5692 13694 5704
rect 14093 5695 14151 5701
rect 14093 5692 14105 5695
rect 13688 5664 14105 5692
rect 13688 5652 13694 5664
rect 14093 5661 14105 5664
rect 14139 5661 14151 5695
rect 14093 5655 14151 5661
rect 18785 5695 18843 5701
rect 18785 5661 18797 5695
rect 18831 5692 18843 5695
rect 18877 5695 18935 5701
rect 18877 5692 18889 5695
rect 18831 5664 18889 5692
rect 18831 5661 18843 5664
rect 18785 5655 18843 5661
rect 18877 5661 18889 5664
rect 18923 5661 18935 5695
rect 18877 5655 18935 5661
rect 21545 5695 21603 5701
rect 21545 5661 21557 5695
rect 21591 5692 21603 5695
rect 21637 5695 21695 5701
rect 21637 5692 21649 5695
rect 21591 5664 21649 5692
rect 21591 5661 21603 5664
rect 21545 5655 21603 5661
rect 21637 5661 21649 5664
rect 21683 5661 21695 5695
rect 21637 5655 21695 5661
rect 28353 5695 28411 5701
rect 28353 5661 28365 5695
rect 28399 5692 28411 5695
rect 31726 5692 31754 5800
rect 34514 5788 34520 5800
rect 34572 5788 34578 5840
rect 38378 5788 38384 5840
rect 38436 5788 38442 5840
rect 36170 5760 36176 5772
rect 34440 5732 36176 5760
rect 34440 5701 34468 5732
rect 36170 5720 36176 5732
rect 36228 5720 36234 5772
rect 28399 5664 31754 5692
rect 34425 5695 34483 5701
rect 28399 5661 28411 5664
rect 28353 5655 28411 5661
rect 34425 5661 34437 5695
rect 34471 5661 34483 5695
rect 34425 5655 34483 5661
rect 35713 5695 35771 5701
rect 35713 5661 35725 5695
rect 35759 5692 35771 5695
rect 36446 5692 36452 5704
rect 35759 5664 36452 5692
rect 35759 5661 35771 5664
rect 35713 5655 35771 5661
rect 36446 5652 36452 5664
rect 36504 5652 36510 5704
rect 36722 5652 36728 5704
rect 36780 5692 36786 5704
rect 36909 5695 36967 5701
rect 36909 5692 36921 5695
rect 36780 5664 36921 5692
rect 36780 5652 36786 5664
rect 36909 5661 36921 5664
rect 36955 5661 36967 5695
rect 36909 5655 36967 5661
rect 36998 5652 37004 5704
rect 37056 5652 37062 5704
rect 37826 5652 37832 5704
rect 37884 5652 37890 5704
rect 38197 5695 38255 5701
rect 38197 5661 38209 5695
rect 38243 5661 38255 5695
rect 38197 5655 38255 5661
rect 11238 5624 11244 5636
rect 4764 5596 7328 5624
rect 7392 5596 11244 5624
rect 4764 5584 4770 5596
rect 6181 5559 6239 5565
rect 6181 5525 6193 5559
rect 6227 5556 6239 5559
rect 7392 5556 7420 5596
rect 11238 5584 11244 5596
rect 11296 5584 11302 5636
rect 12710 5624 12716 5636
rect 12406 5596 12716 5624
rect 6227 5528 7420 5556
rect 7469 5559 7527 5565
rect 6227 5525 6239 5528
rect 6181 5519 6239 5525
rect 7469 5525 7481 5559
rect 7515 5556 7527 5559
rect 12406 5556 12434 5596
rect 12710 5584 12716 5596
rect 12768 5584 12774 5636
rect 16574 5584 16580 5636
rect 16632 5624 16638 5636
rect 20438 5624 20444 5636
rect 16632 5596 20444 5624
rect 16632 5584 16638 5596
rect 20438 5584 20444 5596
rect 20496 5584 20502 5636
rect 38212 5624 38240 5655
rect 22066 5596 38240 5624
rect 7515 5528 12434 5556
rect 7515 5525 7527 5528
rect 7469 5519 7527 5525
rect 13078 5516 13084 5568
rect 13136 5516 13142 5568
rect 13354 5516 13360 5568
rect 13412 5516 13418 5568
rect 13725 5559 13783 5565
rect 13725 5525 13737 5559
rect 13771 5556 13783 5559
rect 21542 5556 21548 5568
rect 13771 5528 21548 5556
rect 13771 5525 13783 5528
rect 13725 5519 13783 5525
rect 21542 5516 21548 5528
rect 21600 5516 21606 5568
rect 21821 5559 21879 5565
rect 21821 5525 21833 5559
rect 21867 5556 21879 5559
rect 22066 5556 22094 5596
rect 21867 5528 22094 5556
rect 21867 5525 21879 5528
rect 21821 5519 21879 5525
rect 38010 5516 38016 5568
rect 38068 5516 38074 5568
rect 1104 5466 38824 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 9010 5466
rect 9062 5414 9074 5466
rect 9126 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 15010 5466
rect 15062 5414 15074 5466
rect 15126 5414 15138 5466
rect 15190 5414 15202 5466
rect 15254 5414 15266 5466
rect 15318 5414 21010 5466
rect 21062 5414 21074 5466
rect 21126 5414 21138 5466
rect 21190 5414 21202 5466
rect 21254 5414 21266 5466
rect 21318 5414 27010 5466
rect 27062 5414 27074 5466
rect 27126 5414 27138 5466
rect 27190 5414 27202 5466
rect 27254 5414 27266 5466
rect 27318 5414 33010 5466
rect 33062 5414 33074 5466
rect 33126 5414 33138 5466
rect 33190 5414 33202 5466
rect 33254 5414 33266 5466
rect 33318 5414 38824 5466
rect 1104 5392 38824 5414
rect 4341 5355 4399 5361
rect 4341 5321 4353 5355
rect 4387 5321 4399 5355
rect 4341 5315 4399 5321
rect 4356 5284 4384 5315
rect 4430 5312 4436 5364
rect 4488 5352 4494 5364
rect 17310 5352 17316 5364
rect 4488 5324 17316 5352
rect 4488 5312 4494 5324
rect 17310 5312 17316 5324
rect 17368 5312 17374 5364
rect 17402 5312 17408 5364
rect 17460 5312 17466 5364
rect 17770 5312 17776 5364
rect 17828 5312 17834 5364
rect 20165 5355 20223 5361
rect 20165 5321 20177 5355
rect 20211 5352 20223 5355
rect 20346 5352 20352 5364
rect 20211 5324 20352 5352
rect 20211 5321 20223 5324
rect 20165 5315 20223 5321
rect 20346 5312 20352 5324
rect 20404 5312 20410 5364
rect 23661 5355 23719 5361
rect 23661 5321 23673 5355
rect 23707 5352 23719 5355
rect 31110 5352 31116 5364
rect 23707 5324 31116 5352
rect 23707 5321 23719 5324
rect 23661 5315 23719 5321
rect 31110 5312 31116 5324
rect 31168 5312 31174 5364
rect 31294 5312 31300 5364
rect 31352 5352 31358 5364
rect 32861 5355 32919 5361
rect 32861 5352 32873 5355
rect 31352 5324 32873 5352
rect 31352 5312 31358 5324
rect 32861 5321 32873 5324
rect 32907 5321 32919 5355
rect 32861 5315 32919 5321
rect 38378 5312 38384 5364
rect 38436 5312 38442 5364
rect 11146 5284 11152 5296
rect 4356 5256 11152 5284
rect 11146 5244 11152 5256
rect 11204 5244 11210 5296
rect 12434 5244 12440 5296
rect 12492 5284 12498 5296
rect 12492 5256 14596 5284
rect 12492 5244 12498 5256
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5185 4215 5219
rect 4157 5179 4215 5185
rect 4433 5219 4491 5225
rect 4433 5185 4445 5219
rect 4479 5185 4491 5219
rect 4433 5179 4491 5185
rect 4709 5219 4767 5225
rect 4709 5185 4721 5219
rect 4755 5216 4767 5219
rect 5258 5216 5264 5228
rect 4755 5188 5264 5216
rect 4755 5185 4767 5188
rect 4709 5179 4767 5185
rect 4172 5080 4200 5179
rect 4448 5148 4476 5179
rect 5258 5176 5264 5188
rect 5316 5176 5322 5228
rect 5350 5176 5356 5228
rect 5408 5216 5414 5228
rect 5537 5219 5595 5225
rect 5537 5216 5549 5219
rect 5408 5188 5549 5216
rect 5408 5176 5414 5188
rect 5537 5185 5549 5188
rect 5583 5185 5595 5219
rect 5537 5179 5595 5185
rect 10502 5176 10508 5228
rect 10560 5216 10566 5228
rect 14568 5225 14596 5256
rect 20530 5244 20536 5296
rect 20588 5284 20594 5296
rect 20588 5256 37872 5284
rect 20588 5244 20594 5256
rect 13725 5219 13783 5225
rect 13725 5216 13737 5219
rect 10560 5188 13737 5216
rect 10560 5176 10566 5188
rect 13725 5185 13737 5188
rect 13771 5185 13783 5219
rect 13725 5179 13783 5185
rect 14001 5219 14059 5225
rect 14001 5185 14013 5219
rect 14047 5185 14059 5219
rect 14001 5179 14059 5185
rect 14277 5219 14335 5225
rect 14277 5185 14289 5219
rect 14323 5185 14335 5219
rect 14277 5179 14335 5185
rect 14553 5219 14611 5225
rect 14553 5185 14565 5219
rect 14599 5185 14611 5219
rect 14553 5179 14611 5185
rect 17497 5219 17555 5225
rect 17497 5185 17509 5219
rect 17543 5216 17555 5219
rect 17589 5219 17647 5225
rect 17589 5216 17601 5219
rect 17543 5188 17601 5216
rect 17543 5185 17555 5188
rect 17497 5179 17555 5185
rect 17589 5185 17601 5188
rect 17635 5185 17647 5219
rect 17589 5179 17647 5185
rect 5810 5148 5816 5160
rect 4448 5120 5816 5148
rect 5810 5108 5816 5120
rect 5868 5108 5874 5160
rect 12158 5108 12164 5160
rect 12216 5148 12222 5160
rect 14016 5148 14044 5179
rect 12216 5120 14044 5148
rect 12216 5108 12222 5120
rect 5534 5080 5540 5092
rect 4172 5052 5540 5080
rect 5534 5040 5540 5052
rect 5592 5040 5598 5092
rect 7558 5080 7564 5092
rect 5644 5052 7564 5080
rect 4614 4972 4620 5024
rect 4672 4972 4678 5024
rect 4893 5015 4951 5021
rect 4893 4981 4905 5015
rect 4939 5012 4951 5015
rect 5644 5012 5672 5052
rect 7558 5040 7564 5052
rect 7616 5040 7622 5092
rect 10226 5040 10232 5092
rect 10284 5080 10290 5092
rect 14292 5080 14320 5179
rect 17770 5176 17776 5228
rect 17828 5216 17834 5228
rect 19797 5219 19855 5225
rect 19797 5216 19809 5219
rect 17828 5188 19809 5216
rect 17828 5176 17834 5188
rect 19797 5185 19809 5188
rect 19843 5216 19855 5219
rect 19981 5219 20039 5225
rect 19981 5216 19993 5219
rect 19843 5188 19993 5216
rect 19843 5185 19855 5188
rect 19797 5179 19855 5185
rect 19981 5185 19993 5188
rect 20027 5185 20039 5219
rect 19981 5179 20039 5185
rect 22925 5219 22983 5225
rect 22925 5185 22937 5219
rect 22971 5216 22983 5219
rect 23017 5219 23075 5225
rect 23017 5216 23029 5219
rect 22971 5188 23029 5216
rect 22971 5185 22983 5188
rect 22925 5179 22983 5185
rect 23017 5185 23029 5188
rect 23063 5185 23075 5219
rect 23017 5179 23075 5185
rect 23385 5219 23443 5225
rect 23385 5185 23397 5219
rect 23431 5216 23443 5219
rect 23477 5219 23535 5225
rect 23477 5216 23489 5219
rect 23431 5188 23489 5216
rect 23431 5185 23443 5188
rect 23385 5179 23443 5185
rect 23477 5185 23489 5188
rect 23523 5185 23535 5219
rect 23477 5179 23535 5185
rect 33045 5219 33103 5225
rect 33045 5185 33057 5219
rect 33091 5216 33103 5219
rect 35986 5216 35992 5228
rect 33091 5188 35992 5216
rect 33091 5185 33103 5188
rect 33045 5179 33103 5185
rect 35986 5176 35992 5188
rect 36044 5176 36050 5228
rect 37844 5225 37872 5256
rect 37829 5219 37887 5225
rect 37829 5185 37841 5219
rect 37875 5185 37887 5219
rect 37829 5179 37887 5185
rect 38197 5219 38255 5225
rect 38197 5185 38209 5219
rect 38243 5185 38255 5219
rect 38197 5179 38255 5185
rect 24854 5148 24860 5160
rect 14476 5120 24860 5148
rect 14476 5089 14504 5120
rect 24854 5108 24860 5120
rect 24912 5108 24918 5160
rect 27890 5108 27896 5160
rect 27948 5148 27954 5160
rect 31386 5148 31392 5160
rect 27948 5120 31392 5148
rect 27948 5108 27954 5120
rect 31386 5108 31392 5120
rect 31444 5108 31450 5160
rect 10284 5052 14320 5080
rect 14461 5083 14519 5089
rect 10284 5040 10290 5052
rect 14461 5049 14473 5083
rect 14507 5049 14519 5083
rect 14461 5043 14519 5049
rect 19610 5040 19616 5092
rect 19668 5080 19674 5092
rect 38212 5080 38240 5179
rect 19668 5052 38240 5080
rect 19668 5040 19674 5052
rect 4939 4984 5672 5012
rect 4939 4981 4951 4984
rect 4893 4975 4951 4981
rect 5718 4972 5724 5024
rect 5776 4972 5782 5024
rect 13814 4972 13820 5024
rect 13872 5012 13878 5024
rect 13909 5015 13967 5021
rect 13909 5012 13921 5015
rect 13872 4984 13921 5012
rect 13872 4972 13878 4984
rect 13909 4981 13921 4984
rect 13955 4981 13967 5015
rect 13909 4975 13967 4981
rect 14185 5015 14243 5021
rect 14185 4981 14197 5015
rect 14231 5012 14243 5015
rect 14366 5012 14372 5024
rect 14231 4984 14372 5012
rect 14231 4981 14243 4984
rect 14185 4975 14243 4981
rect 14366 4972 14372 4984
rect 14424 4972 14430 5024
rect 14737 5015 14795 5021
rect 14737 4981 14749 5015
rect 14783 5012 14795 5015
rect 17586 5012 17592 5024
rect 14783 4984 17592 5012
rect 14783 4981 14795 4984
rect 14737 4975 14795 4981
rect 17586 4972 17592 4984
rect 17644 4972 17650 5024
rect 22830 4972 22836 5024
rect 22888 4972 22894 5024
rect 23198 4972 23204 5024
rect 23256 4972 23262 5024
rect 23290 4972 23296 5024
rect 23348 4972 23354 5024
rect 28166 4972 28172 5024
rect 28224 5012 28230 5024
rect 30558 5012 30564 5024
rect 28224 4984 30564 5012
rect 28224 4972 28230 4984
rect 30558 4972 30564 4984
rect 30616 4972 30622 5024
rect 38013 5015 38071 5021
rect 38013 4981 38025 5015
rect 38059 5012 38071 5015
rect 39114 5012 39120 5024
rect 38059 4984 39120 5012
rect 38059 4981 38071 4984
rect 38013 4975 38071 4981
rect 39114 4972 39120 4984
rect 39172 4972 39178 5024
rect 1104 4922 38824 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 13950 4922
rect 14002 4870 14014 4922
rect 14066 4870 14078 4922
rect 14130 4870 14142 4922
rect 14194 4870 14206 4922
rect 14258 4870 19950 4922
rect 20002 4870 20014 4922
rect 20066 4870 20078 4922
rect 20130 4870 20142 4922
rect 20194 4870 20206 4922
rect 20258 4870 25950 4922
rect 26002 4870 26014 4922
rect 26066 4870 26078 4922
rect 26130 4870 26142 4922
rect 26194 4870 26206 4922
rect 26258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 37950 4922
rect 38002 4870 38014 4922
rect 38066 4870 38078 4922
rect 38130 4870 38142 4922
rect 38194 4870 38206 4922
rect 38258 4870 38824 4922
rect 1104 4848 38824 4870
rect 4430 4768 4436 4820
rect 4488 4768 4494 4820
rect 4614 4768 4620 4820
rect 4672 4808 4678 4820
rect 11514 4808 11520 4820
rect 4672 4780 11520 4808
rect 4672 4768 4678 4780
rect 11514 4768 11520 4780
rect 11572 4768 11578 4820
rect 15470 4768 15476 4820
rect 15528 4768 15534 4820
rect 17862 4768 17868 4820
rect 17920 4808 17926 4820
rect 19337 4811 19395 4817
rect 19337 4808 19349 4811
rect 17920 4780 19349 4808
rect 17920 4768 17926 4780
rect 19337 4777 19349 4780
rect 19383 4777 19395 4811
rect 19337 4771 19395 4777
rect 19610 4768 19616 4820
rect 19668 4768 19674 4820
rect 27522 4808 27528 4820
rect 22066 4780 27528 4808
rect 2774 4700 2780 4752
rect 2832 4740 2838 4752
rect 5350 4740 5356 4752
rect 2832 4712 5356 4740
rect 2832 4700 2838 4712
rect 5350 4700 5356 4712
rect 5408 4700 5414 4752
rect 11054 4700 11060 4752
rect 11112 4740 11118 4752
rect 21634 4740 21640 4752
rect 11112 4712 21640 4740
rect 11112 4700 11118 4712
rect 21634 4700 21640 4712
rect 21692 4700 21698 4752
rect 21729 4743 21787 4749
rect 21729 4709 21741 4743
rect 21775 4740 21787 4743
rect 22066 4740 22094 4780
rect 27522 4768 27528 4780
rect 27580 4768 27586 4820
rect 27614 4768 27620 4820
rect 27672 4808 27678 4820
rect 29549 4811 29607 4817
rect 29549 4808 29561 4811
rect 27672 4780 29561 4808
rect 27672 4768 27678 4780
rect 29549 4777 29561 4780
rect 29595 4777 29607 4811
rect 29549 4771 29607 4777
rect 30742 4768 30748 4820
rect 30800 4768 30806 4820
rect 30834 4768 30840 4820
rect 30892 4808 30898 4820
rect 35342 4808 35348 4820
rect 30892 4780 35348 4808
rect 30892 4768 30898 4780
rect 35342 4768 35348 4780
rect 35400 4768 35406 4820
rect 25498 4740 25504 4752
rect 21775 4712 22094 4740
rect 22388 4712 25504 4740
rect 21775 4709 21787 4712
rect 21729 4703 21787 4709
rect 13814 4632 13820 4684
rect 13872 4672 13878 4684
rect 22388 4672 22416 4712
rect 25498 4700 25504 4712
rect 25556 4700 25562 4752
rect 26326 4700 26332 4752
rect 26384 4740 26390 4752
rect 28261 4743 28319 4749
rect 28261 4740 28273 4743
rect 26384 4712 28273 4740
rect 26384 4700 26390 4712
rect 28261 4709 28273 4712
rect 28307 4709 28319 4743
rect 28261 4703 28319 4709
rect 31110 4700 31116 4752
rect 31168 4740 31174 4752
rect 38194 4740 38200 4752
rect 31168 4712 38200 4740
rect 31168 4700 31174 4712
rect 38194 4700 38200 4712
rect 38252 4700 38258 4752
rect 38378 4700 38384 4752
rect 38436 4700 38442 4752
rect 13872 4644 19564 4672
rect 13872 4632 13878 4644
rect 2866 4564 2872 4616
rect 2924 4604 2930 4616
rect 4249 4607 4307 4613
rect 4249 4604 4261 4607
rect 2924 4576 4261 4604
rect 2924 4564 2930 4576
rect 4249 4573 4261 4576
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 9674 4564 9680 4616
rect 9732 4604 9738 4616
rect 15013 4607 15071 4613
rect 15013 4604 15025 4607
rect 9732 4576 15025 4604
rect 9732 4564 9738 4576
rect 15013 4573 15025 4576
rect 15059 4573 15071 4607
rect 15013 4567 15071 4573
rect 15289 4607 15347 4613
rect 15289 4573 15301 4607
rect 15335 4604 15347 4607
rect 15562 4604 15568 4616
rect 15335 4576 15568 4604
rect 15335 4573 15347 4576
rect 15289 4567 15347 4573
rect 15562 4564 15568 4576
rect 15620 4564 15626 4616
rect 19337 4607 19395 4613
rect 19337 4573 19349 4607
rect 19383 4604 19395 4607
rect 19429 4607 19487 4613
rect 19429 4604 19441 4607
rect 19383 4576 19441 4604
rect 19383 4573 19395 4576
rect 19337 4567 19395 4573
rect 19429 4573 19441 4576
rect 19475 4573 19487 4607
rect 19536 4604 19564 4644
rect 19720 4644 22416 4672
rect 19720 4604 19748 4644
rect 23198 4632 23204 4684
rect 23256 4672 23262 4684
rect 35618 4672 35624 4684
rect 23256 4644 29132 4672
rect 23256 4632 23262 4644
rect 19536 4576 19748 4604
rect 19429 4567 19487 4573
rect 21358 4564 21364 4616
rect 21416 4604 21422 4616
rect 21545 4607 21603 4613
rect 21545 4604 21557 4607
rect 21416 4576 21557 4604
rect 21416 4564 21422 4576
rect 21545 4573 21557 4576
rect 21591 4573 21603 4607
rect 21545 4567 21603 4573
rect 23569 4607 23627 4613
rect 23569 4573 23581 4607
rect 23615 4573 23627 4607
rect 25682 4604 25688 4616
rect 23569 4567 23627 4573
rect 23676 4576 25688 4604
rect 5718 4496 5724 4548
rect 5776 4536 5782 4548
rect 13814 4536 13820 4548
rect 5776 4508 13820 4536
rect 5776 4496 5782 4508
rect 13814 4496 13820 4508
rect 13872 4496 13878 4548
rect 15470 4496 15476 4548
rect 15528 4536 15534 4548
rect 15528 4508 19288 4536
rect 15528 4496 15534 4508
rect 15197 4471 15255 4477
rect 15197 4437 15209 4471
rect 15243 4468 15255 4471
rect 17862 4468 17868 4480
rect 15243 4440 17868 4468
rect 15243 4437 15255 4440
rect 15197 4431 15255 4437
rect 17862 4428 17868 4440
rect 17920 4428 17926 4480
rect 19260 4468 19288 4508
rect 21634 4496 21640 4548
rect 21692 4536 21698 4548
rect 23477 4539 23535 4545
rect 23477 4536 23489 4539
rect 21692 4508 23489 4536
rect 21692 4496 21698 4508
rect 23477 4505 23489 4508
rect 23523 4536 23535 4539
rect 23584 4536 23612 4567
rect 23523 4508 23612 4536
rect 23523 4505 23535 4508
rect 23477 4499 23535 4505
rect 23676 4468 23704 4576
rect 25682 4564 25688 4576
rect 25740 4564 25746 4616
rect 27985 4607 28043 4613
rect 27709 4583 27767 4589
rect 27709 4580 27721 4583
rect 27632 4552 27721 4580
rect 19260 4440 23704 4468
rect 23750 4428 23756 4480
rect 23808 4428 23814 4480
rect 24210 4428 24216 4480
rect 24268 4468 24274 4480
rect 27632 4477 27660 4552
rect 27709 4549 27721 4552
rect 27755 4549 27767 4583
rect 27985 4573 27997 4607
rect 28031 4604 28043 4607
rect 28261 4607 28319 4613
rect 28261 4604 28273 4607
rect 28031 4576 28273 4604
rect 28031 4573 28043 4576
rect 27985 4567 28043 4573
rect 28261 4573 28273 4576
rect 28307 4573 28319 4607
rect 28261 4567 28319 4573
rect 28994 4564 29000 4616
rect 29052 4564 29058 4616
rect 27709 4543 27767 4549
rect 27798 4496 27804 4548
rect 27856 4536 27862 4548
rect 29104 4536 29132 4644
rect 30944 4644 35624 4672
rect 29733 4607 29791 4613
rect 29733 4573 29745 4607
rect 29779 4604 29791 4607
rect 30834 4604 30840 4616
rect 29779 4576 30840 4604
rect 29779 4573 29791 4576
rect 29733 4567 29791 4573
rect 30834 4564 30840 4576
rect 30892 4564 30898 4616
rect 30944 4613 30972 4644
rect 35618 4632 35624 4644
rect 35676 4632 35682 4684
rect 30929 4607 30987 4613
rect 30929 4573 30941 4607
rect 30975 4573 30987 4607
rect 37829 4607 37887 4613
rect 37829 4604 37841 4607
rect 30929 4567 30987 4573
rect 31036 4576 37841 4604
rect 31036 4536 31064 4576
rect 37829 4573 37841 4576
rect 37875 4573 37887 4607
rect 37829 4567 37887 4573
rect 38197 4607 38255 4613
rect 38197 4573 38209 4607
rect 38243 4573 38255 4607
rect 38197 4567 38255 4573
rect 38212 4536 38240 4567
rect 27856 4508 28948 4536
rect 29104 4508 31064 4536
rect 31726 4508 38240 4536
rect 27856 4496 27862 4508
rect 27617 4471 27675 4477
rect 27617 4468 27629 4471
rect 24268 4440 27629 4468
rect 24268 4428 24274 4440
rect 27617 4437 27629 4440
rect 27663 4437 27675 4471
rect 27617 4431 27675 4437
rect 27890 4428 27896 4480
rect 27948 4428 27954 4480
rect 28166 4428 28172 4480
rect 28224 4428 28230 4480
rect 28810 4428 28816 4480
rect 28868 4428 28874 4480
rect 28920 4468 28948 4508
rect 31726 4468 31754 4508
rect 28920 4440 31754 4468
rect 38010 4428 38016 4480
rect 38068 4428 38074 4480
rect 1104 4378 38824 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 9010 4378
rect 9062 4326 9074 4378
rect 9126 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 15010 4378
rect 15062 4326 15074 4378
rect 15126 4326 15138 4378
rect 15190 4326 15202 4378
rect 15254 4326 15266 4378
rect 15318 4326 21010 4378
rect 21062 4326 21074 4378
rect 21126 4326 21138 4378
rect 21190 4326 21202 4378
rect 21254 4326 21266 4378
rect 21318 4326 27010 4378
rect 27062 4326 27074 4378
rect 27126 4326 27138 4378
rect 27190 4326 27202 4378
rect 27254 4326 27266 4378
rect 27318 4326 33010 4378
rect 33062 4326 33074 4378
rect 33126 4326 33138 4378
rect 33190 4326 33202 4378
rect 33254 4326 33266 4378
rect 33318 4326 38824 4378
rect 1104 4304 38824 4326
rect 566 4224 572 4276
rect 624 4264 630 4276
rect 19426 4264 19432 4276
rect 624 4236 19432 4264
rect 624 4224 630 4236
rect 19426 4224 19432 4236
rect 19484 4224 19490 4276
rect 19610 4224 19616 4276
rect 19668 4264 19674 4276
rect 19668 4236 23704 4264
rect 19668 4224 19674 4236
rect 5718 4156 5724 4208
rect 5776 4196 5782 4208
rect 15838 4196 15844 4208
rect 5776 4168 15844 4196
rect 5776 4156 5782 4168
rect 15838 4156 15844 4168
rect 15896 4156 15902 4208
rect 19794 4156 19800 4208
rect 19852 4196 19858 4208
rect 22370 4196 22376 4208
rect 19852 4168 22376 4196
rect 19852 4156 19858 4168
rect 22370 4156 22376 4168
rect 22428 4156 22434 4208
rect 23676 4196 23704 4236
rect 23750 4224 23756 4276
rect 23808 4264 23814 4276
rect 23808 4236 37872 4264
rect 23808 4224 23814 4236
rect 24394 4196 24400 4208
rect 23676 4168 24400 4196
rect 24394 4156 24400 4168
rect 24452 4156 24458 4208
rect 28994 4156 29000 4208
rect 29052 4196 29058 4208
rect 29638 4196 29644 4208
rect 29052 4168 29644 4196
rect 29052 4156 29058 4168
rect 29638 4156 29644 4168
rect 29696 4156 29702 4208
rect 2869 4131 2927 4137
rect 2869 4097 2881 4131
rect 2915 4128 2927 4131
rect 3602 4128 3608 4140
rect 2915 4100 3608 4128
rect 2915 4097 2927 4100
rect 2869 4091 2927 4097
rect 3602 4088 3608 4100
rect 3660 4088 3666 4140
rect 9398 4088 9404 4140
rect 9456 4128 9462 4140
rect 15933 4131 15991 4137
rect 15933 4128 15945 4131
rect 9456 4100 15945 4128
rect 9456 4088 9462 4100
rect 15933 4097 15945 4100
rect 15979 4097 15991 4131
rect 15933 4091 15991 4097
rect 19153 4131 19211 4137
rect 19153 4097 19165 4131
rect 19199 4128 19211 4131
rect 19245 4131 19303 4137
rect 19245 4128 19257 4131
rect 19199 4100 19257 4128
rect 19199 4097 19211 4100
rect 19153 4091 19211 4097
rect 19245 4097 19257 4100
rect 19291 4097 19303 4131
rect 19245 4091 19303 4097
rect 20714 4088 20720 4140
rect 20772 4128 20778 4140
rect 21821 4131 21879 4137
rect 21821 4128 21833 4131
rect 20772 4100 21833 4128
rect 20772 4088 20778 4100
rect 21821 4097 21833 4100
rect 21867 4128 21879 4131
rect 22097 4131 22155 4137
rect 22097 4128 22109 4131
rect 21867 4100 22109 4128
rect 21867 4097 21879 4100
rect 21821 4091 21879 4097
rect 22097 4097 22109 4100
rect 22143 4097 22155 4131
rect 22097 4091 22155 4097
rect 25593 4131 25651 4137
rect 25593 4097 25605 4131
rect 25639 4128 25651 4131
rect 25685 4131 25743 4137
rect 25685 4128 25697 4131
rect 25639 4100 25697 4128
rect 25639 4097 25651 4100
rect 25593 4091 25651 4097
rect 25685 4097 25697 4100
rect 25731 4097 25743 4131
rect 25685 4091 25743 4097
rect 26421 4131 26479 4137
rect 26421 4097 26433 4131
rect 26467 4128 26479 4131
rect 26513 4131 26571 4137
rect 26513 4128 26525 4131
rect 26467 4100 26525 4128
rect 26467 4097 26479 4100
rect 26421 4091 26479 4097
rect 26513 4097 26525 4100
rect 26559 4097 26571 4131
rect 26513 4091 26571 4097
rect 27065 4131 27123 4137
rect 27065 4097 27077 4131
rect 27111 4097 27123 4131
rect 27065 4091 27123 4097
rect 27709 4131 27767 4137
rect 27709 4097 27721 4131
rect 27755 4128 27767 4131
rect 27798 4128 27804 4140
rect 27755 4100 27804 4128
rect 27755 4097 27767 4100
rect 27709 4091 27767 4097
rect 7650 4020 7656 4072
rect 7708 4060 7714 4072
rect 19061 4063 19119 4069
rect 19061 4060 19073 4063
rect 7708 4032 19073 4060
rect 7708 4020 7714 4032
rect 19061 4029 19073 4032
rect 19107 4029 19119 4063
rect 19061 4023 19119 4029
rect 19334 4020 19340 4072
rect 19392 4060 19398 4072
rect 23842 4060 23848 4072
rect 19392 4032 23848 4060
rect 19392 4020 19398 4032
rect 23842 4020 23848 4032
rect 23900 4020 23906 4072
rect 24946 4020 24952 4072
rect 25004 4060 25010 4072
rect 27080 4060 27108 4091
rect 27798 4088 27804 4100
rect 27856 4088 27862 4140
rect 28261 4131 28319 4137
rect 28261 4097 28273 4131
rect 28307 4097 28319 4131
rect 28261 4091 28319 4097
rect 25004 4032 27108 4060
rect 28276 4060 28304 4091
rect 28350 4088 28356 4140
rect 28408 4088 28414 4140
rect 28813 4131 28871 4137
rect 28813 4097 28825 4131
rect 28859 4128 28871 4131
rect 29089 4131 29147 4137
rect 29089 4128 29101 4131
rect 28859 4100 29101 4128
rect 28859 4097 28871 4100
rect 28813 4091 28871 4097
rect 29089 4097 29101 4100
rect 29135 4097 29147 4131
rect 29089 4091 29147 4097
rect 29178 4088 29184 4140
rect 29236 4128 29242 4140
rect 37844 4137 37872 4236
rect 29457 4131 29515 4137
rect 29457 4128 29469 4131
rect 29236 4100 29469 4128
rect 29236 4088 29242 4100
rect 29457 4097 29469 4100
rect 29503 4097 29515 4131
rect 29457 4091 29515 4097
rect 29733 4131 29791 4137
rect 29733 4097 29745 4131
rect 29779 4128 29791 4131
rect 29825 4131 29883 4137
rect 29825 4128 29837 4131
rect 29779 4100 29837 4128
rect 29779 4097 29791 4100
rect 29733 4091 29791 4097
rect 29825 4097 29837 4100
rect 29871 4097 29883 4131
rect 29825 4091 29883 4097
rect 30193 4131 30251 4137
rect 30193 4097 30205 4131
rect 30239 4128 30251 4131
rect 30469 4131 30527 4137
rect 30469 4128 30481 4131
rect 30239 4100 30481 4128
rect 30239 4097 30251 4100
rect 30193 4091 30251 4097
rect 30469 4097 30481 4100
rect 30515 4097 30527 4131
rect 30469 4091 30527 4097
rect 30745 4131 30803 4137
rect 30745 4097 30757 4131
rect 30791 4128 30803 4131
rect 30837 4131 30895 4137
rect 30837 4128 30849 4131
rect 30791 4100 30849 4128
rect 30791 4097 30803 4100
rect 30745 4091 30803 4097
rect 30837 4097 30849 4100
rect 30883 4097 30895 4131
rect 30837 4091 30895 4097
rect 31205 4131 31263 4137
rect 31205 4097 31217 4131
rect 31251 4097 31263 4131
rect 31205 4091 31263 4097
rect 37829 4131 37887 4137
rect 37829 4097 37841 4131
rect 37875 4097 37887 4131
rect 37829 4091 37887 4097
rect 28534 4060 28540 4072
rect 28276 4032 28540 4060
rect 25004 4020 25010 4032
rect 28534 4020 28540 4032
rect 28592 4020 28598 4072
rect 29546 4020 29552 4072
rect 29604 4060 29610 4072
rect 30101 4063 30159 4069
rect 30101 4060 30113 4063
rect 29604 4032 30113 4060
rect 29604 4020 29610 4032
rect 30101 4029 30113 4032
rect 30147 4029 30159 4063
rect 30101 4023 30159 4029
rect 30282 4020 30288 4072
rect 30340 4060 30346 4072
rect 31220 4060 31248 4091
rect 38194 4088 38200 4140
rect 38252 4088 38258 4140
rect 30340 4032 31248 4060
rect 30340 4020 30346 4032
rect 31294 4020 31300 4072
rect 31352 4060 31358 4072
rect 37458 4060 37464 4072
rect 31352 4032 37464 4060
rect 31352 4020 31358 4032
rect 37458 4020 37464 4032
rect 37516 4020 37522 4072
rect 16117 3995 16175 4001
rect 16117 3961 16129 3995
rect 16163 3992 16175 3995
rect 16163 3964 21956 3992
rect 16163 3961 16175 3964
rect 16117 3955 16175 3961
rect 3050 3884 3056 3936
rect 3108 3884 3114 3936
rect 5626 3884 5632 3936
rect 5684 3924 5690 3936
rect 19334 3924 19340 3936
rect 5684 3896 19340 3924
rect 5684 3884 5690 3896
rect 19334 3884 19340 3896
rect 19392 3884 19398 3936
rect 19429 3927 19487 3933
rect 19429 3893 19441 3927
rect 19475 3924 19487 3927
rect 20530 3924 20536 3936
rect 19475 3896 20536 3924
rect 19475 3893 19487 3896
rect 19429 3887 19487 3893
rect 20530 3884 20536 3896
rect 20588 3884 20594 3936
rect 21928 3924 21956 3964
rect 22002 3952 22008 4004
rect 22060 3952 22066 4004
rect 23474 3952 23480 4004
rect 23532 3992 23538 4004
rect 25406 3992 25412 4004
rect 23532 3964 25412 3992
rect 23532 3952 23538 3964
rect 25406 3952 25412 3964
rect 25464 3952 25470 4004
rect 25774 3952 25780 4004
rect 25832 3992 25838 4004
rect 28077 3995 28135 4001
rect 28077 3992 28089 3995
rect 25832 3964 28089 3992
rect 25832 3952 25838 3964
rect 28077 3961 28089 3964
rect 28123 3961 28135 3995
rect 28077 3955 28135 3961
rect 28258 3952 28264 4004
rect 28316 3992 28322 4004
rect 28721 3995 28779 4001
rect 28721 3992 28733 3995
rect 28316 3964 28733 3992
rect 28316 3952 28322 3964
rect 28721 3961 28733 3964
rect 28767 3961 28779 3995
rect 28721 3955 28779 3961
rect 29365 3995 29423 4001
rect 29365 3961 29377 3995
rect 29411 3992 29423 3995
rect 30466 3992 30472 4004
rect 29411 3964 30472 3992
rect 29411 3961 29423 3964
rect 29365 3955 29423 3961
rect 30466 3952 30472 3964
rect 30524 3952 30530 4004
rect 38378 3952 38384 4004
rect 38436 3952 38442 4004
rect 23198 3924 23204 3936
rect 21928 3896 23204 3924
rect 23198 3884 23204 3896
rect 23256 3884 23262 3936
rect 25038 3884 25044 3936
rect 25096 3924 25102 3936
rect 25501 3927 25559 3933
rect 25501 3924 25513 3927
rect 25096 3896 25513 3924
rect 25096 3884 25102 3896
rect 25501 3893 25513 3896
rect 25547 3893 25559 3927
rect 25501 3887 25559 3893
rect 25866 3884 25872 3936
rect 25924 3884 25930 3936
rect 26418 3884 26424 3936
rect 26476 3884 26482 3936
rect 26694 3884 26700 3936
rect 26752 3884 26758 3936
rect 27249 3927 27307 3933
rect 27249 3893 27261 3927
rect 27295 3924 27307 3927
rect 27430 3924 27436 3936
rect 27295 3896 27436 3924
rect 27295 3893 27307 3896
rect 27249 3887 27307 3893
rect 27430 3884 27436 3896
rect 27488 3884 27494 3936
rect 27890 3884 27896 3936
rect 27948 3884 27954 3936
rect 28537 3927 28595 3933
rect 28537 3893 28549 3927
rect 28583 3924 28595 3927
rect 28626 3924 28632 3936
rect 28583 3896 28632 3924
rect 28583 3893 28595 3896
rect 28537 3887 28595 3893
rect 28626 3884 28632 3896
rect 28684 3884 28690 3936
rect 28810 3884 28816 3936
rect 28868 3924 28874 3936
rect 28905 3927 28963 3933
rect 28905 3924 28917 3927
rect 28868 3896 28917 3924
rect 28868 3884 28874 3896
rect 28905 3893 28917 3896
rect 28951 3893 28963 3927
rect 28905 3887 28963 3893
rect 29454 3884 29460 3936
rect 29512 3924 29518 3936
rect 29641 3927 29699 3933
rect 29641 3924 29653 3927
rect 29512 3896 29653 3924
rect 29512 3884 29518 3896
rect 29641 3893 29653 3896
rect 29687 3893 29699 3927
rect 29641 3887 29699 3893
rect 30006 3884 30012 3936
rect 30064 3884 30070 3936
rect 30190 3884 30196 3936
rect 30248 3924 30254 3936
rect 30285 3927 30343 3933
rect 30285 3924 30297 3927
rect 30248 3896 30297 3924
rect 30248 3884 30254 3896
rect 30285 3893 30297 3896
rect 30331 3893 30343 3927
rect 30285 3887 30343 3893
rect 30374 3884 30380 3936
rect 30432 3924 30438 3936
rect 30561 3927 30619 3933
rect 30561 3924 30573 3927
rect 30432 3896 30573 3924
rect 30432 3884 30438 3896
rect 30561 3893 30573 3896
rect 30607 3893 30619 3927
rect 30561 3887 30619 3893
rect 30834 3884 30840 3936
rect 30892 3884 30898 3936
rect 31021 3927 31079 3933
rect 31021 3893 31033 3927
rect 31067 3924 31079 3927
rect 31110 3924 31116 3936
rect 31067 3896 31116 3924
rect 31067 3893 31079 3896
rect 31021 3887 31079 3893
rect 31110 3884 31116 3896
rect 31168 3884 31174 3936
rect 38013 3927 38071 3933
rect 38013 3893 38025 3927
rect 38059 3924 38071 3927
rect 39114 3924 39120 3936
rect 38059 3896 39120 3924
rect 38059 3893 38071 3896
rect 38013 3887 38071 3893
rect 39114 3884 39120 3896
rect 39172 3884 39178 3936
rect 1104 3834 38824 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 13950 3834
rect 14002 3782 14014 3834
rect 14066 3782 14078 3834
rect 14130 3782 14142 3834
rect 14194 3782 14206 3834
rect 14258 3782 19950 3834
rect 20002 3782 20014 3834
rect 20066 3782 20078 3834
rect 20130 3782 20142 3834
rect 20194 3782 20206 3834
rect 20258 3782 25950 3834
rect 26002 3782 26014 3834
rect 26066 3782 26078 3834
rect 26130 3782 26142 3834
rect 26194 3782 26206 3834
rect 26258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 37950 3834
rect 38002 3782 38014 3834
rect 38066 3782 38078 3834
rect 38130 3782 38142 3834
rect 38194 3782 38206 3834
rect 38258 3782 38824 3834
rect 1104 3760 38824 3782
rect 17037 3723 17095 3729
rect 17037 3689 17049 3723
rect 17083 3720 17095 3723
rect 23474 3720 23480 3732
rect 17083 3692 23480 3720
rect 17083 3689 17095 3692
rect 17037 3683 17095 3689
rect 23474 3680 23480 3692
rect 23532 3680 23538 3732
rect 23658 3680 23664 3732
rect 23716 3720 23722 3732
rect 24857 3723 24915 3729
rect 24857 3720 24869 3723
rect 23716 3692 24869 3720
rect 23716 3680 23722 3692
rect 24857 3689 24869 3692
rect 24903 3689 24915 3723
rect 24857 3683 24915 3689
rect 25866 3680 25872 3732
rect 25924 3720 25930 3732
rect 28626 3720 28632 3732
rect 25924 3692 28632 3720
rect 25924 3680 25930 3692
rect 28626 3680 28632 3692
rect 28684 3680 28690 3732
rect 28718 3680 28724 3732
rect 28776 3720 28782 3732
rect 31018 3720 31024 3732
rect 28776 3692 31024 3720
rect 28776 3680 28782 3692
rect 31018 3680 31024 3692
rect 31076 3680 31082 3732
rect 3050 3612 3056 3664
rect 3108 3652 3114 3664
rect 15378 3652 15384 3664
rect 3108 3624 15384 3652
rect 3108 3612 3114 3624
rect 15378 3612 15384 3624
rect 15436 3612 15442 3664
rect 16577 3655 16635 3661
rect 16577 3621 16589 3655
rect 16623 3621 16635 3655
rect 16577 3615 16635 3621
rect 17681 3655 17739 3661
rect 17681 3621 17693 3655
rect 17727 3652 17739 3655
rect 20346 3652 20352 3664
rect 17727 3624 20352 3652
rect 17727 3621 17739 3624
rect 17681 3615 17739 3621
rect 16592 3584 16620 3615
rect 20346 3612 20352 3624
rect 20404 3612 20410 3664
rect 20714 3612 20720 3664
rect 20772 3652 20778 3664
rect 21726 3652 21732 3664
rect 20772 3624 21732 3652
rect 20772 3612 20778 3624
rect 21726 3612 21732 3624
rect 21784 3612 21790 3664
rect 21818 3612 21824 3664
rect 21876 3612 21882 3664
rect 23569 3655 23627 3661
rect 23569 3621 23581 3655
rect 23615 3621 23627 3655
rect 23569 3615 23627 3621
rect 23845 3655 23903 3661
rect 23845 3621 23857 3655
rect 23891 3652 23903 3655
rect 23891 3624 31754 3652
rect 23891 3621 23903 3624
rect 23845 3615 23903 3621
rect 23474 3584 23480 3596
rect 16592 3556 23480 3584
rect 23474 3544 23480 3556
rect 23532 3544 23538 3596
rect 23584 3584 23612 3615
rect 23584 3556 29868 3584
rect 3418 3476 3424 3528
rect 3476 3516 3482 3528
rect 3789 3519 3847 3525
rect 3789 3516 3801 3519
rect 3476 3488 3801 3516
rect 3476 3476 3482 3488
rect 3789 3485 3801 3488
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 8846 3476 8852 3528
rect 8904 3516 8910 3528
rect 16393 3519 16451 3525
rect 16393 3516 16405 3519
rect 8904 3488 16405 3516
rect 8904 3476 8910 3488
rect 16393 3485 16405 3488
rect 16439 3485 16451 3519
rect 16393 3479 16451 3485
rect 16850 3476 16856 3528
rect 16908 3476 16914 3528
rect 16942 3476 16948 3528
rect 17000 3516 17006 3528
rect 17497 3519 17555 3525
rect 17497 3516 17509 3519
rect 17000 3488 17509 3516
rect 17000 3476 17006 3488
rect 17497 3485 17509 3488
rect 17543 3485 17555 3519
rect 17497 3479 17555 3485
rect 17770 3476 17776 3528
rect 17828 3476 17834 3528
rect 19334 3476 19340 3528
rect 19392 3516 19398 3528
rect 20714 3516 20720 3528
rect 19392 3488 20720 3516
rect 19392 3476 19398 3488
rect 20714 3476 20720 3488
rect 20772 3476 20778 3528
rect 20993 3519 21051 3525
rect 20993 3485 21005 3519
rect 21039 3516 21051 3519
rect 21085 3519 21143 3525
rect 21085 3516 21097 3519
rect 21039 3488 21097 3516
rect 21039 3485 21051 3488
rect 20993 3479 21051 3485
rect 21085 3485 21097 3488
rect 21131 3485 21143 3519
rect 21085 3479 21143 3485
rect 21634 3476 21640 3528
rect 21692 3476 21698 3528
rect 21726 3476 21732 3528
rect 21784 3516 21790 3528
rect 22097 3519 22155 3525
rect 22097 3516 22109 3519
rect 21784 3488 22109 3516
rect 21784 3476 21790 3488
rect 22097 3485 22109 3488
rect 22143 3485 22155 3519
rect 22097 3479 22155 3485
rect 22557 3519 22615 3525
rect 22557 3485 22569 3519
rect 22603 3516 22615 3519
rect 22649 3519 22707 3525
rect 22649 3516 22661 3519
rect 22603 3488 22661 3516
rect 22603 3485 22615 3488
rect 22557 3479 22615 3485
rect 22649 3485 22661 3488
rect 22695 3485 22707 3519
rect 22649 3479 22707 3485
rect 23109 3519 23167 3525
rect 23109 3485 23121 3519
rect 23155 3516 23167 3519
rect 23385 3519 23443 3525
rect 23385 3516 23397 3519
rect 23155 3488 23397 3516
rect 23155 3485 23167 3488
rect 23109 3479 23167 3485
rect 23385 3485 23397 3488
rect 23431 3485 23443 3519
rect 23385 3479 23443 3485
rect 23658 3476 23664 3528
rect 23716 3476 23722 3528
rect 23937 3519 23995 3525
rect 23937 3485 23949 3519
rect 23983 3485 23995 3519
rect 23937 3479 23995 3485
rect 9582 3408 9588 3460
rect 9640 3448 9646 3460
rect 22465 3451 22523 3457
rect 22465 3448 22477 3451
rect 9640 3420 22477 3448
rect 9640 3408 9646 3420
rect 22465 3417 22477 3420
rect 22511 3417 22523 3451
rect 22465 3411 22523 3417
rect 23293 3451 23351 3457
rect 23293 3417 23305 3451
rect 23339 3448 23351 3451
rect 23952 3448 23980 3479
rect 24394 3476 24400 3528
rect 24452 3516 24458 3528
rect 24673 3519 24731 3525
rect 24673 3516 24685 3519
rect 24452 3488 24685 3516
rect 24452 3476 24458 3488
rect 24673 3485 24685 3488
rect 24719 3485 24731 3519
rect 24673 3479 24731 3485
rect 28813 3519 28871 3525
rect 28813 3485 28825 3519
rect 28859 3516 28871 3519
rect 29089 3519 29147 3525
rect 29089 3516 29101 3519
rect 28859 3488 29101 3516
rect 28859 3485 28871 3488
rect 28813 3479 28871 3485
rect 29089 3485 29101 3488
rect 29135 3485 29147 3519
rect 29089 3479 29147 3485
rect 29270 3476 29276 3528
rect 29328 3516 29334 3528
rect 29733 3519 29791 3525
rect 29733 3516 29745 3519
rect 29328 3488 29745 3516
rect 29328 3476 29334 3488
rect 29733 3485 29745 3488
rect 29779 3485 29791 3519
rect 29733 3479 29791 3485
rect 29638 3448 29644 3460
rect 23339 3420 23980 3448
rect 24136 3420 29644 3448
rect 23339 3417 23351 3420
rect 23293 3411 23351 3417
rect 3970 3340 3976 3392
rect 4028 3340 4034 3392
rect 12618 3340 12624 3392
rect 12676 3380 12682 3392
rect 17678 3380 17684 3392
rect 12676 3352 17684 3380
rect 12676 3340 12682 3352
rect 17678 3340 17684 3352
rect 17736 3340 17742 3392
rect 17954 3340 17960 3392
rect 18012 3340 18018 3392
rect 20622 3340 20628 3392
rect 20680 3380 20686 3392
rect 20901 3383 20959 3389
rect 20901 3380 20913 3383
rect 20680 3352 20913 3380
rect 20680 3340 20686 3352
rect 20901 3349 20913 3352
rect 20947 3349 20959 3383
rect 20901 3343 20959 3349
rect 21269 3383 21327 3389
rect 21269 3349 21281 3383
rect 21315 3380 21327 3383
rect 21726 3380 21732 3392
rect 21315 3352 21732 3380
rect 21315 3349 21327 3352
rect 21269 3343 21327 3349
rect 21726 3340 21732 3352
rect 21784 3340 21790 3392
rect 22281 3383 22339 3389
rect 22281 3349 22293 3383
rect 22327 3380 22339 3383
rect 22738 3380 22744 3392
rect 22327 3352 22744 3380
rect 22327 3349 22339 3352
rect 22281 3343 22339 3349
rect 22738 3340 22744 3352
rect 22796 3340 22802 3392
rect 22830 3340 22836 3392
rect 22888 3340 22894 3392
rect 23014 3340 23020 3392
rect 23072 3340 23078 3392
rect 23106 3340 23112 3392
rect 23164 3380 23170 3392
rect 24136 3389 24164 3420
rect 29638 3408 29644 3420
rect 29696 3408 29702 3460
rect 29840 3448 29868 3556
rect 30009 3519 30067 3525
rect 30009 3485 30021 3519
rect 30055 3516 30067 3519
rect 30101 3519 30159 3525
rect 30101 3516 30113 3519
rect 30055 3488 30113 3516
rect 30055 3485 30067 3488
rect 30009 3479 30067 3485
rect 30101 3485 30113 3488
rect 30147 3485 30159 3519
rect 31726 3516 31754 3624
rect 38378 3612 38384 3664
rect 38436 3612 38442 3664
rect 35894 3544 35900 3596
rect 35952 3584 35958 3596
rect 35952 3556 38240 3584
rect 35952 3544 35958 3556
rect 38212 3525 38240 3556
rect 37829 3519 37887 3525
rect 37829 3516 37841 3519
rect 31726 3488 37841 3516
rect 30101 3479 30159 3485
rect 37829 3485 37841 3488
rect 37875 3485 37887 3519
rect 37829 3479 37887 3485
rect 38197 3519 38255 3525
rect 38197 3485 38209 3519
rect 38243 3485 38255 3519
rect 38197 3479 38255 3485
rect 37918 3448 37924 3460
rect 29840 3420 37924 3448
rect 37918 3408 37924 3420
rect 37976 3408 37982 3460
rect 23201 3383 23259 3389
rect 23201 3380 23213 3383
rect 23164 3352 23213 3380
rect 23164 3340 23170 3352
rect 23201 3349 23213 3352
rect 23247 3349 23259 3383
rect 23201 3343 23259 3349
rect 24121 3383 24179 3389
rect 24121 3349 24133 3383
rect 24167 3349 24179 3383
rect 24121 3343 24179 3349
rect 24486 3340 24492 3392
rect 24544 3380 24550 3392
rect 24581 3383 24639 3389
rect 24581 3380 24593 3383
rect 24544 3352 24593 3380
rect 24544 3340 24550 3352
rect 24581 3349 24593 3352
rect 24627 3349 24639 3383
rect 24581 3343 24639 3349
rect 25314 3340 25320 3392
rect 25372 3380 25378 3392
rect 28721 3383 28779 3389
rect 28721 3380 28733 3383
rect 25372 3352 28733 3380
rect 25372 3340 25378 3352
rect 28721 3349 28733 3352
rect 28767 3349 28779 3383
rect 28721 3343 28779 3349
rect 28902 3340 28908 3392
rect 28960 3340 28966 3392
rect 29546 3340 29552 3392
rect 29604 3340 29610 3392
rect 29822 3340 29828 3392
rect 29880 3340 29886 3392
rect 30193 3383 30251 3389
rect 30193 3349 30205 3383
rect 30239 3380 30251 3383
rect 30282 3380 30288 3392
rect 30239 3352 30288 3380
rect 30239 3349 30251 3352
rect 30193 3343 30251 3349
rect 30282 3340 30288 3352
rect 30340 3340 30346 3392
rect 38010 3340 38016 3392
rect 38068 3340 38074 3392
rect 1104 3290 38824 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 9010 3290
rect 9062 3238 9074 3290
rect 9126 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 15010 3290
rect 15062 3238 15074 3290
rect 15126 3238 15138 3290
rect 15190 3238 15202 3290
rect 15254 3238 15266 3290
rect 15318 3238 21010 3290
rect 21062 3238 21074 3290
rect 21126 3238 21138 3290
rect 21190 3238 21202 3290
rect 21254 3238 21266 3290
rect 21318 3238 27010 3290
rect 27062 3238 27074 3290
rect 27126 3238 27138 3290
rect 27190 3238 27202 3290
rect 27254 3238 27266 3290
rect 27318 3238 33010 3290
rect 33062 3238 33074 3290
rect 33126 3238 33138 3290
rect 33190 3238 33202 3290
rect 33254 3238 33266 3290
rect 33318 3238 38824 3290
rect 1104 3216 38824 3238
rect 10962 3136 10968 3188
rect 11020 3176 11026 3188
rect 21634 3176 21640 3188
rect 11020 3148 21640 3176
rect 11020 3136 11026 3148
rect 21634 3136 21640 3148
rect 21692 3136 21698 3188
rect 22557 3179 22615 3185
rect 22557 3145 22569 3179
rect 22603 3176 22615 3179
rect 23290 3176 23296 3188
rect 22603 3148 23296 3176
rect 22603 3145 22615 3148
rect 22557 3139 22615 3145
rect 23290 3136 23296 3148
rect 23348 3136 23354 3188
rect 27062 3176 27068 3188
rect 23400 3148 27068 3176
rect 8294 3068 8300 3120
rect 8352 3108 8358 3120
rect 16942 3108 16948 3120
rect 8352 3080 16948 3108
rect 8352 3068 8358 3080
rect 16942 3068 16948 3080
rect 17000 3068 17006 3120
rect 17770 3108 17776 3120
rect 17052 3080 17776 3108
rect 8570 3000 8576 3052
rect 8628 3040 8634 3052
rect 17052 3040 17080 3080
rect 17770 3068 17776 3080
rect 17828 3068 17834 3120
rect 17954 3068 17960 3120
rect 18012 3108 18018 3120
rect 23400 3108 23428 3148
rect 27062 3136 27068 3148
rect 27120 3136 27126 3188
rect 29546 3176 29552 3188
rect 28828 3148 29552 3176
rect 18012 3080 23428 3108
rect 18012 3068 18018 3080
rect 23474 3068 23480 3120
rect 23532 3108 23538 3120
rect 23532 3080 26188 3108
rect 23532 3068 23538 3080
rect 8628 3012 17080 3040
rect 17497 3043 17555 3049
rect 8628 3000 8634 3012
rect 17497 3009 17509 3043
rect 17543 3009 17555 3043
rect 17497 3003 17555 3009
rect 10778 2932 10784 2984
rect 10836 2972 10842 2984
rect 13630 2972 13636 2984
rect 10836 2944 13636 2972
rect 10836 2932 10842 2944
rect 13630 2932 13636 2944
rect 13688 2932 13694 2984
rect 3970 2864 3976 2916
rect 4028 2904 4034 2916
rect 17512 2904 17540 3003
rect 18598 3000 18604 3052
rect 18656 3000 18662 3052
rect 19429 3043 19487 3049
rect 19429 3009 19441 3043
rect 19475 3040 19487 3043
rect 19702 3040 19708 3052
rect 19475 3012 19708 3040
rect 19475 3009 19487 3012
rect 19429 3003 19487 3009
rect 19702 3000 19708 3012
rect 19760 3000 19766 3052
rect 20732 3012 22232 3040
rect 17678 2932 17684 2984
rect 17736 2972 17742 2984
rect 19242 2972 19248 2984
rect 17736 2944 19248 2972
rect 17736 2932 17742 2944
rect 19242 2932 19248 2944
rect 19300 2932 19306 2984
rect 4028 2876 17540 2904
rect 4028 2864 4034 2876
rect 17586 2864 17592 2916
rect 17644 2904 17650 2916
rect 20732 2904 20760 3012
rect 21542 2932 21548 2984
rect 21600 2972 21606 2984
rect 22204 2972 22232 3012
rect 22370 3000 22376 3052
rect 22428 3000 22434 3052
rect 22741 3043 22799 3049
rect 22741 3040 22753 3043
rect 22480 3012 22753 3040
rect 22480 2972 22508 3012
rect 22741 3009 22753 3012
rect 22787 3009 22799 3043
rect 23293 3043 23351 3049
rect 23293 3040 23305 3043
rect 22741 3003 22799 3009
rect 22848 3012 23305 3040
rect 22848 2972 22876 3012
rect 23293 3009 23305 3012
rect 23339 3009 23351 3043
rect 23293 3003 23351 3009
rect 23842 3000 23848 3052
rect 23900 3000 23906 3052
rect 24854 3000 24860 3052
rect 24912 3040 24918 3052
rect 26160 3049 26188 3080
rect 24949 3043 25007 3049
rect 24949 3040 24961 3043
rect 24912 3012 24961 3040
rect 24912 3000 24918 3012
rect 24949 3009 24961 3012
rect 24995 3009 25007 3043
rect 25777 3043 25835 3049
rect 25777 3040 25789 3043
rect 24949 3003 25007 3009
rect 25056 3012 25789 3040
rect 21600 2944 22140 2972
rect 22204 2944 22508 2972
rect 22572 2944 22876 2972
rect 21600 2932 21606 2944
rect 17644 2876 20760 2904
rect 22112 2904 22140 2944
rect 22572 2904 22600 2944
rect 23198 2932 23204 2984
rect 23256 2972 23262 2984
rect 25056 2972 25084 3012
rect 25777 3009 25789 3012
rect 25823 3009 25835 3043
rect 25777 3003 25835 3009
rect 26145 3043 26203 3049
rect 26145 3009 26157 3043
rect 26191 3009 26203 3043
rect 26145 3003 26203 3009
rect 27430 3000 27436 3052
rect 27488 3000 27494 3052
rect 28537 3043 28595 3049
rect 28537 3009 28549 3043
rect 28583 3040 28595 3043
rect 28828 3040 28856 3148
rect 29546 3136 29552 3148
rect 29604 3136 29610 3188
rect 29638 3136 29644 3188
rect 29696 3176 29702 3188
rect 29696 3148 37872 3176
rect 29696 3136 29702 3148
rect 29822 3108 29828 3120
rect 28920 3080 29828 3108
rect 28920 3049 28948 3080
rect 29822 3068 29828 3080
rect 29880 3068 29886 3120
rect 28583 3012 28856 3040
rect 28905 3043 28963 3049
rect 28583 3009 28595 3012
rect 28537 3003 28595 3009
rect 28905 3009 28917 3043
rect 28951 3009 28963 3043
rect 28905 3003 28963 3009
rect 29641 3043 29699 3049
rect 29641 3009 29653 3043
rect 29687 3040 29699 3043
rect 30374 3040 30380 3052
rect 29687 3012 30380 3040
rect 29687 3009 29699 3012
rect 29641 3003 29699 3009
rect 30374 3000 30380 3012
rect 30432 3000 30438 3052
rect 30469 3043 30527 3049
rect 30469 3009 30481 3043
rect 30515 3040 30527 3043
rect 30558 3040 30564 3052
rect 30515 3012 30564 3040
rect 30515 3009 30527 3012
rect 30469 3003 30527 3009
rect 30558 3000 30564 3012
rect 30616 3000 30622 3052
rect 31021 3043 31079 3049
rect 31021 3009 31033 3043
rect 31067 3009 31079 3043
rect 31021 3003 31079 3009
rect 23256 2944 25084 2972
rect 25792 2944 26464 2972
rect 23256 2932 23262 2944
rect 22112 2876 22600 2904
rect 17644 2864 17650 2876
rect 22830 2864 22836 2916
rect 22888 2904 22894 2916
rect 25792 2904 25820 2944
rect 22888 2876 25820 2904
rect 22888 2864 22894 2876
rect 25866 2864 25872 2916
rect 25924 2904 25930 2916
rect 26329 2907 26387 2913
rect 26329 2904 26341 2907
rect 25924 2876 26341 2904
rect 25924 2864 25930 2876
rect 26329 2873 26341 2876
rect 26375 2873 26387 2907
rect 26436 2904 26464 2944
rect 26694 2932 26700 2984
rect 26752 2972 26758 2984
rect 31036 2972 31064 3003
rect 37458 3000 37464 3052
rect 37516 3000 37522 3052
rect 37844 3049 37872 3148
rect 38378 3136 38384 3188
rect 38436 3136 38442 3188
rect 37829 3043 37887 3049
rect 37829 3009 37841 3043
rect 37875 3009 37887 3043
rect 37829 3003 37887 3009
rect 37918 3000 37924 3052
rect 37976 3040 37982 3052
rect 38197 3043 38255 3049
rect 38197 3040 38209 3043
rect 37976 3012 38209 3040
rect 37976 3000 37982 3012
rect 38197 3009 38209 3012
rect 38243 3009 38255 3043
rect 38197 3003 38255 3009
rect 26752 2944 31064 2972
rect 26752 2932 26758 2944
rect 31294 2904 31300 2916
rect 26436 2876 31300 2904
rect 26329 2867 26387 2873
rect 31294 2864 31300 2876
rect 31352 2864 31358 2916
rect 11238 2796 11244 2848
rect 11296 2836 11302 2848
rect 11606 2836 11612 2848
rect 11296 2808 11612 2836
rect 11296 2796 11302 2808
rect 11606 2796 11612 2808
rect 11664 2796 11670 2848
rect 17402 2796 17408 2848
rect 17460 2836 17466 2848
rect 17681 2839 17739 2845
rect 17681 2836 17693 2839
rect 17460 2808 17693 2836
rect 17460 2796 17466 2808
rect 17681 2805 17693 2808
rect 17727 2805 17739 2839
rect 17681 2799 17739 2805
rect 18506 2796 18512 2848
rect 18564 2836 18570 2848
rect 18785 2839 18843 2845
rect 18785 2836 18797 2839
rect 18564 2808 18797 2836
rect 18564 2796 18570 2808
rect 18785 2805 18797 2808
rect 18831 2805 18843 2839
rect 18785 2799 18843 2805
rect 19334 2796 19340 2848
rect 19392 2836 19398 2848
rect 19613 2839 19671 2845
rect 19613 2836 19625 2839
rect 19392 2808 19625 2836
rect 19392 2796 19398 2808
rect 19613 2805 19625 2808
rect 19659 2805 19671 2839
rect 19613 2799 19671 2805
rect 22646 2796 22652 2848
rect 22704 2836 22710 2848
rect 22925 2839 22983 2845
rect 22925 2836 22937 2839
rect 22704 2808 22937 2836
rect 22704 2796 22710 2808
rect 22925 2805 22937 2808
rect 22971 2805 22983 2839
rect 22925 2799 22983 2805
rect 23198 2796 23204 2848
rect 23256 2836 23262 2848
rect 23477 2839 23535 2845
rect 23477 2836 23489 2839
rect 23256 2808 23489 2836
rect 23256 2796 23262 2808
rect 23477 2805 23489 2808
rect 23523 2805 23535 2839
rect 23477 2799 23535 2805
rect 23750 2796 23756 2848
rect 23808 2836 23814 2848
rect 24029 2839 24087 2845
rect 24029 2836 24041 2839
rect 23808 2808 24041 2836
rect 23808 2796 23814 2808
rect 24029 2805 24041 2808
rect 24075 2805 24087 2839
rect 24029 2799 24087 2805
rect 24854 2796 24860 2848
rect 24912 2836 24918 2848
rect 25133 2839 25191 2845
rect 25133 2836 25145 2839
rect 24912 2808 25145 2836
rect 24912 2796 24918 2808
rect 25133 2805 25145 2808
rect 25179 2805 25191 2839
rect 25133 2799 25191 2805
rect 25682 2796 25688 2848
rect 25740 2836 25746 2848
rect 25961 2839 26019 2845
rect 25961 2836 25973 2839
rect 25740 2808 25973 2836
rect 25740 2796 25746 2808
rect 25961 2805 25973 2808
rect 26007 2805 26019 2839
rect 25961 2799 26019 2805
rect 26878 2796 26884 2848
rect 26936 2836 26942 2848
rect 27249 2839 27307 2845
rect 27249 2836 27261 2839
rect 26936 2808 27261 2836
rect 26936 2796 26942 2808
rect 27249 2805 27261 2808
rect 27295 2805 27307 2839
rect 27249 2799 27307 2805
rect 28166 2796 28172 2848
rect 28224 2836 28230 2848
rect 28353 2839 28411 2845
rect 28353 2836 28365 2839
rect 28224 2808 28365 2836
rect 28224 2796 28230 2808
rect 28353 2805 28365 2808
rect 28399 2805 28411 2839
rect 28353 2799 28411 2805
rect 28442 2796 28448 2848
rect 28500 2836 28506 2848
rect 28721 2839 28779 2845
rect 28721 2836 28733 2839
rect 28500 2808 28733 2836
rect 28500 2796 28506 2808
rect 28721 2805 28733 2808
rect 28767 2805 28779 2839
rect 28721 2799 28779 2805
rect 29270 2796 29276 2848
rect 29328 2836 29334 2848
rect 29457 2839 29515 2845
rect 29457 2836 29469 2839
rect 29328 2808 29469 2836
rect 29328 2796 29334 2808
rect 29457 2805 29469 2808
rect 29503 2805 29515 2839
rect 29457 2799 29515 2805
rect 30374 2796 30380 2848
rect 30432 2836 30438 2848
rect 30653 2839 30711 2845
rect 30653 2836 30665 2839
rect 30432 2808 30665 2836
rect 30432 2796 30438 2808
rect 30653 2805 30665 2808
rect 30699 2805 30711 2839
rect 30653 2799 30711 2805
rect 30926 2796 30932 2848
rect 30984 2836 30990 2848
rect 31205 2839 31263 2845
rect 31205 2836 31217 2839
rect 30984 2808 31217 2836
rect 30984 2796 30990 2808
rect 31205 2805 31217 2808
rect 31251 2805 31263 2839
rect 31205 2799 31263 2805
rect 37645 2839 37703 2845
rect 37645 2805 37657 2839
rect 37691 2836 37703 2839
rect 37826 2836 37832 2848
rect 37691 2808 37832 2836
rect 37691 2805 37703 2808
rect 37645 2799 37703 2805
rect 37826 2796 37832 2808
rect 37884 2796 37890 2848
rect 38013 2839 38071 2845
rect 38013 2805 38025 2839
rect 38059 2836 38071 2839
rect 39114 2836 39120 2848
rect 38059 2808 39120 2836
rect 38059 2805 38071 2808
rect 38013 2799 38071 2805
rect 39114 2796 39120 2808
rect 39172 2796 39178 2848
rect 1104 2746 38824 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 13950 2746
rect 14002 2694 14014 2746
rect 14066 2694 14078 2746
rect 14130 2694 14142 2746
rect 14194 2694 14206 2746
rect 14258 2694 19950 2746
rect 20002 2694 20014 2746
rect 20066 2694 20078 2746
rect 20130 2694 20142 2746
rect 20194 2694 20206 2746
rect 20258 2694 25950 2746
rect 26002 2694 26014 2746
rect 26066 2694 26078 2746
rect 26130 2694 26142 2746
rect 26194 2694 26206 2746
rect 26258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 37950 2746
rect 38002 2694 38014 2746
rect 38066 2694 38078 2746
rect 38130 2694 38142 2746
rect 38194 2694 38206 2746
rect 38258 2694 38824 2746
rect 1104 2672 38824 2694
rect 14274 2592 14280 2644
rect 14332 2632 14338 2644
rect 14332 2604 20852 2632
rect 14332 2592 14338 2604
rect 7558 2524 7564 2576
rect 7616 2564 7622 2576
rect 7616 2536 18460 2564
rect 7616 2524 7622 2536
rect 9490 2456 9496 2508
rect 9548 2496 9554 2508
rect 9548 2468 18368 2496
rect 9548 2456 9554 2468
rect 15378 2388 15384 2440
rect 15436 2428 15442 2440
rect 16945 2431 17003 2437
rect 16945 2428 16957 2431
rect 15436 2400 16957 2428
rect 15436 2388 15442 2400
rect 16945 2397 16957 2400
rect 16991 2397 17003 2431
rect 16945 2391 17003 2397
rect 17310 2388 17316 2440
rect 17368 2388 17374 2440
rect 17681 2431 17739 2437
rect 17681 2397 17693 2431
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 13814 2320 13820 2372
rect 13872 2360 13878 2372
rect 17696 2360 17724 2391
rect 18046 2388 18052 2440
rect 18104 2388 18110 2440
rect 13872 2332 17724 2360
rect 18340 2360 18368 2468
rect 18432 2437 18460 2536
rect 18874 2524 18880 2576
rect 18932 2564 18938 2576
rect 19610 2564 19616 2576
rect 18932 2536 19616 2564
rect 18932 2524 18938 2536
rect 19610 2524 19616 2536
rect 19668 2524 19674 2576
rect 18598 2456 18604 2508
rect 18656 2496 18662 2508
rect 20824 2496 20852 2604
rect 21818 2592 21824 2644
rect 21876 2632 21882 2644
rect 22462 2632 22468 2644
rect 21876 2604 22468 2632
rect 21876 2592 21882 2604
rect 22462 2592 22468 2604
rect 22520 2592 22526 2644
rect 22756 2604 23244 2632
rect 21542 2524 21548 2576
rect 21600 2564 21606 2576
rect 22373 2567 22431 2573
rect 22373 2564 22385 2567
rect 21600 2536 22385 2564
rect 21600 2524 21606 2536
rect 22373 2533 22385 2536
rect 22419 2533 22431 2567
rect 22373 2527 22431 2533
rect 22756 2496 22784 2604
rect 23109 2567 23167 2573
rect 23109 2564 23121 2567
rect 18656 2468 19748 2496
rect 20824 2468 22784 2496
rect 22848 2536 23121 2564
rect 18656 2456 18662 2468
rect 18417 2431 18475 2437
rect 18417 2397 18429 2431
rect 18463 2397 18475 2431
rect 18417 2391 18475 2397
rect 18782 2388 18788 2440
rect 18840 2388 18846 2440
rect 19242 2388 19248 2440
rect 19300 2388 19306 2440
rect 19610 2388 19616 2440
rect 19668 2388 19674 2440
rect 19720 2428 19748 2468
rect 19981 2431 20039 2437
rect 19981 2428 19993 2431
rect 19720 2400 19993 2428
rect 19981 2397 19993 2400
rect 20027 2397 20039 2431
rect 19981 2391 20039 2397
rect 20349 2431 20407 2437
rect 20349 2397 20361 2431
rect 20395 2428 20407 2431
rect 20438 2428 20444 2440
rect 20395 2400 20444 2428
rect 20395 2397 20407 2400
rect 20349 2391 20407 2397
rect 20438 2388 20444 2400
rect 20496 2388 20502 2440
rect 20530 2388 20536 2440
rect 20588 2428 20594 2440
rect 20717 2431 20775 2437
rect 20717 2428 20729 2431
rect 20588 2400 20729 2428
rect 20588 2388 20594 2400
rect 20717 2397 20729 2400
rect 20763 2397 20775 2431
rect 20717 2391 20775 2397
rect 20806 2388 20812 2440
rect 20864 2428 20870 2440
rect 21085 2431 21143 2437
rect 21085 2428 21097 2431
rect 20864 2400 21097 2428
rect 20864 2388 20870 2400
rect 21085 2397 21097 2400
rect 21131 2397 21143 2431
rect 21085 2391 21143 2397
rect 21821 2431 21879 2437
rect 21821 2397 21833 2431
rect 21867 2397 21879 2431
rect 21821 2391 21879 2397
rect 21836 2360 21864 2391
rect 22186 2388 22192 2440
rect 22244 2388 22250 2440
rect 22278 2388 22284 2440
rect 22336 2428 22342 2440
rect 22557 2431 22615 2437
rect 22557 2428 22569 2431
rect 22336 2400 22569 2428
rect 22336 2388 22342 2400
rect 22557 2397 22569 2400
rect 22603 2397 22615 2431
rect 22557 2391 22615 2397
rect 18340 2332 21864 2360
rect 13872 2320 13878 2332
rect 22094 2320 22100 2372
rect 22152 2360 22158 2372
rect 22848 2360 22876 2536
rect 23109 2533 23121 2536
rect 23155 2533 23167 2567
rect 23109 2527 23167 2533
rect 23216 2496 23244 2604
rect 23474 2592 23480 2644
rect 23532 2632 23538 2644
rect 24581 2635 24639 2641
rect 24581 2632 24593 2635
rect 23532 2604 24593 2632
rect 23532 2592 23538 2604
rect 24581 2601 24593 2604
rect 24627 2601 24639 2635
rect 24581 2595 24639 2601
rect 24670 2592 24676 2644
rect 24728 2632 24734 2644
rect 25685 2635 25743 2641
rect 25685 2632 25697 2635
rect 24728 2604 25697 2632
rect 24728 2592 24734 2604
rect 25685 2601 25697 2604
rect 25731 2601 25743 2635
rect 25685 2595 25743 2601
rect 26142 2592 26148 2644
rect 26200 2632 26206 2644
rect 26326 2632 26332 2644
rect 26200 2604 26332 2632
rect 26200 2592 26206 2604
rect 26326 2592 26332 2604
rect 26384 2592 26390 2644
rect 26786 2592 26792 2644
rect 26844 2632 26850 2644
rect 27893 2635 27951 2641
rect 27893 2632 27905 2635
rect 26844 2604 27905 2632
rect 26844 2592 26850 2604
rect 27893 2601 27905 2604
rect 27939 2601 27951 2635
rect 27893 2595 27951 2601
rect 27982 2592 27988 2644
rect 28040 2632 28046 2644
rect 28905 2635 28963 2641
rect 28905 2632 28917 2635
rect 28040 2604 28917 2632
rect 28040 2592 28046 2604
rect 28905 2601 28917 2604
rect 28951 2601 28963 2635
rect 28905 2595 28963 2601
rect 29822 2592 29828 2644
rect 29880 2632 29886 2644
rect 30837 2635 30895 2641
rect 30837 2632 30849 2635
rect 29880 2604 30849 2632
rect 29880 2592 29886 2604
rect 30837 2601 30849 2604
rect 30883 2601 30895 2635
rect 30837 2595 30895 2601
rect 24026 2524 24032 2576
rect 24084 2564 24090 2576
rect 24949 2567 25007 2573
rect 24949 2564 24961 2567
rect 24084 2536 24961 2564
rect 24084 2524 24090 2536
rect 24949 2533 24961 2536
rect 24995 2533 25007 2567
rect 24949 2527 25007 2533
rect 25130 2524 25136 2576
rect 25188 2564 25194 2576
rect 26053 2567 26111 2573
rect 26053 2564 26065 2567
rect 25188 2536 26065 2564
rect 25188 2524 25194 2536
rect 26053 2533 26065 2536
rect 26099 2533 26111 2567
rect 26053 2527 26111 2533
rect 26234 2524 26240 2576
rect 26292 2564 26298 2576
rect 27157 2567 27215 2573
rect 27157 2564 27169 2567
rect 26292 2536 27169 2564
rect 26292 2524 26298 2536
rect 27157 2533 27169 2536
rect 27203 2533 27215 2567
rect 27157 2527 27215 2533
rect 27338 2524 27344 2576
rect 27396 2564 27402 2576
rect 28261 2567 28319 2573
rect 28261 2564 28273 2567
rect 27396 2536 28273 2564
rect 27396 2524 27402 2536
rect 28261 2533 28273 2536
rect 28307 2533 28319 2567
rect 28261 2527 28319 2533
rect 28718 2524 28724 2576
rect 28776 2564 28782 2576
rect 29641 2567 29699 2573
rect 29641 2564 29653 2567
rect 28776 2536 29653 2564
rect 28776 2524 28782 2536
rect 29641 2533 29653 2536
rect 29687 2533 29699 2567
rect 29641 2527 29699 2533
rect 30098 2524 30104 2576
rect 30156 2564 30162 2576
rect 30156 2536 30420 2564
rect 30156 2524 30162 2536
rect 23216 2468 25176 2496
rect 22922 2388 22928 2440
rect 22980 2388 22986 2440
rect 23014 2388 23020 2440
rect 23072 2428 23078 2440
rect 23293 2431 23351 2437
rect 23293 2428 23305 2431
rect 23072 2400 23305 2428
rect 23072 2388 23078 2400
rect 23293 2397 23305 2400
rect 23339 2397 23351 2431
rect 23293 2391 23351 2397
rect 23658 2388 23664 2440
rect 23716 2388 23722 2440
rect 24394 2388 24400 2440
rect 24452 2388 24458 2440
rect 24762 2388 24768 2440
rect 24820 2388 24826 2440
rect 25148 2437 25176 2468
rect 25406 2456 25412 2508
rect 25464 2496 25470 2508
rect 25464 2468 27016 2496
rect 25464 2456 25470 2468
rect 25133 2431 25191 2437
rect 25133 2397 25145 2431
rect 25179 2397 25191 2431
rect 25133 2391 25191 2397
rect 25498 2388 25504 2440
rect 25556 2388 25562 2440
rect 25774 2388 25780 2440
rect 25832 2428 25838 2440
rect 25869 2431 25927 2437
rect 25869 2428 25881 2431
rect 25832 2400 25881 2428
rect 25832 2388 25838 2400
rect 25869 2397 25881 2400
rect 25915 2397 25927 2431
rect 25869 2391 25927 2397
rect 25958 2388 25964 2440
rect 26016 2428 26022 2440
rect 26988 2437 27016 2468
rect 30006 2456 30012 2508
rect 30064 2496 30070 2508
rect 30392 2496 30420 2536
rect 30466 2524 30472 2576
rect 30524 2524 30530 2576
rect 30650 2524 30656 2576
rect 30708 2564 30714 2576
rect 31573 2567 31631 2573
rect 31573 2564 31585 2567
rect 30708 2536 31585 2564
rect 30708 2524 30714 2536
rect 31573 2533 31585 2536
rect 31619 2533 31631 2567
rect 31573 2527 31631 2533
rect 33502 2524 33508 2576
rect 33560 2564 33566 2576
rect 33560 2536 37872 2564
rect 33560 2524 33566 2536
rect 30064 2468 30328 2496
rect 30392 2468 31248 2496
rect 30064 2456 30070 2468
rect 26237 2431 26295 2437
rect 26237 2428 26249 2431
rect 26016 2400 26249 2428
rect 26016 2388 26022 2400
rect 26237 2397 26249 2400
rect 26283 2397 26295 2431
rect 26237 2391 26295 2397
rect 26973 2431 27031 2437
rect 26973 2397 26985 2431
rect 27019 2397 27031 2431
rect 26973 2391 27031 2397
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27341 2431 27399 2437
rect 27341 2428 27353 2431
rect 27120 2400 27353 2428
rect 27120 2388 27126 2400
rect 27341 2397 27353 2400
rect 27387 2397 27399 2431
rect 27341 2391 27399 2397
rect 27706 2388 27712 2440
rect 27764 2388 27770 2440
rect 27890 2388 27896 2440
rect 27948 2428 27954 2440
rect 28077 2431 28135 2437
rect 28077 2428 28089 2431
rect 27948 2400 28089 2428
rect 27948 2388 27954 2400
rect 28077 2397 28089 2400
rect 28123 2397 28135 2431
rect 28077 2391 28135 2397
rect 28721 2431 28779 2437
rect 28721 2397 28733 2431
rect 28767 2428 28779 2431
rect 28810 2428 28816 2440
rect 28767 2400 28816 2428
rect 28767 2397 28779 2400
rect 28721 2391 28779 2397
rect 28810 2388 28816 2400
rect 28868 2388 28874 2440
rect 28902 2388 28908 2440
rect 28960 2428 28966 2440
rect 29089 2431 29147 2437
rect 29089 2428 29101 2431
rect 28960 2400 29101 2428
rect 28960 2388 28966 2400
rect 29089 2397 29101 2400
rect 29135 2397 29147 2431
rect 29089 2391 29147 2397
rect 29825 2431 29883 2437
rect 29825 2397 29837 2431
rect 29871 2428 29883 2431
rect 29871 2400 30144 2428
rect 29871 2397 29883 2400
rect 29825 2391 29883 2397
rect 22152 2332 22876 2360
rect 22940 2332 23888 2360
rect 22152 2320 22158 2332
rect 22940 2304 22968 2332
rect 17126 2252 17132 2304
rect 17184 2252 17190 2304
rect 17497 2295 17555 2301
rect 17497 2261 17509 2295
rect 17543 2292 17555 2295
rect 17678 2292 17684 2304
rect 17543 2264 17684 2292
rect 17543 2261 17555 2264
rect 17497 2255 17555 2261
rect 17678 2252 17684 2264
rect 17736 2252 17742 2304
rect 17865 2295 17923 2301
rect 17865 2261 17877 2295
rect 17911 2292 17923 2295
rect 17954 2292 17960 2304
rect 17911 2264 17960 2292
rect 17911 2261 17923 2264
rect 17865 2255 17923 2261
rect 17954 2252 17960 2264
rect 18012 2252 18018 2304
rect 18230 2252 18236 2304
rect 18288 2252 18294 2304
rect 18601 2295 18659 2301
rect 18601 2261 18613 2295
rect 18647 2292 18659 2295
rect 18782 2292 18788 2304
rect 18647 2264 18788 2292
rect 18647 2261 18659 2264
rect 18601 2255 18659 2261
rect 18782 2252 18788 2264
rect 18840 2252 18846 2304
rect 18969 2295 19027 2301
rect 18969 2261 18981 2295
rect 19015 2292 19027 2295
rect 19058 2292 19064 2304
rect 19015 2264 19064 2292
rect 19015 2261 19027 2264
rect 18969 2255 19027 2261
rect 19058 2252 19064 2264
rect 19116 2252 19122 2304
rect 19429 2295 19487 2301
rect 19429 2261 19441 2295
rect 19475 2292 19487 2295
rect 19610 2292 19616 2304
rect 19475 2264 19616 2292
rect 19475 2261 19487 2264
rect 19429 2255 19487 2261
rect 19610 2252 19616 2264
rect 19668 2252 19674 2304
rect 19797 2295 19855 2301
rect 19797 2261 19809 2295
rect 19843 2292 19855 2295
rect 19886 2292 19892 2304
rect 19843 2264 19892 2292
rect 19843 2261 19855 2264
rect 19797 2255 19855 2261
rect 19886 2252 19892 2264
rect 19944 2252 19950 2304
rect 20162 2252 20168 2304
rect 20220 2252 20226 2304
rect 20438 2252 20444 2304
rect 20496 2292 20502 2304
rect 20533 2295 20591 2301
rect 20533 2292 20545 2295
rect 20496 2264 20545 2292
rect 20496 2252 20502 2264
rect 20533 2261 20545 2264
rect 20579 2261 20591 2295
rect 20533 2255 20591 2261
rect 20714 2252 20720 2304
rect 20772 2292 20778 2304
rect 20901 2295 20959 2301
rect 20901 2292 20913 2295
rect 20772 2264 20913 2292
rect 20772 2252 20778 2264
rect 20901 2261 20913 2264
rect 20947 2261 20959 2295
rect 20901 2255 20959 2261
rect 20990 2252 20996 2304
rect 21048 2292 21054 2304
rect 21269 2295 21327 2301
rect 21269 2292 21281 2295
rect 21048 2264 21281 2292
rect 21048 2252 21054 2264
rect 21269 2261 21281 2264
rect 21315 2261 21327 2295
rect 21269 2255 21327 2261
rect 21358 2252 21364 2304
rect 21416 2292 21422 2304
rect 22005 2295 22063 2301
rect 22005 2292 22017 2295
rect 21416 2264 22017 2292
rect 21416 2252 21422 2264
rect 22005 2261 22017 2264
rect 22051 2261 22063 2295
rect 22005 2255 22063 2261
rect 22462 2252 22468 2304
rect 22520 2292 22526 2304
rect 22741 2295 22799 2301
rect 22741 2292 22753 2295
rect 22520 2264 22753 2292
rect 22520 2252 22526 2264
rect 22741 2261 22753 2264
rect 22787 2261 22799 2295
rect 22741 2255 22799 2261
rect 22922 2252 22928 2304
rect 22980 2252 22986 2304
rect 23014 2252 23020 2304
rect 23072 2292 23078 2304
rect 23860 2301 23888 2332
rect 24302 2320 24308 2372
rect 24360 2360 24366 2372
rect 24360 2332 25360 2360
rect 24360 2320 24366 2332
rect 25332 2301 25360 2332
rect 25406 2320 25412 2372
rect 25464 2360 25470 2372
rect 25464 2332 26464 2360
rect 25464 2320 25470 2332
rect 26436 2301 26464 2332
rect 27614 2320 27620 2372
rect 27672 2360 27678 2372
rect 27672 2332 28580 2360
rect 27672 2320 27678 2332
rect 23477 2295 23535 2301
rect 23477 2292 23489 2295
rect 23072 2264 23489 2292
rect 23072 2252 23078 2264
rect 23477 2261 23489 2264
rect 23523 2261 23535 2295
rect 23477 2255 23535 2261
rect 23845 2295 23903 2301
rect 23845 2261 23857 2295
rect 23891 2261 23903 2295
rect 23845 2255 23903 2261
rect 25317 2295 25375 2301
rect 25317 2261 25329 2295
rect 25363 2261 25375 2295
rect 25317 2255 25375 2261
rect 26421 2295 26479 2301
rect 26421 2261 26433 2295
rect 26467 2261 26479 2295
rect 26421 2255 26479 2261
rect 26510 2252 26516 2304
rect 26568 2292 26574 2304
rect 28552 2301 28580 2332
rect 27525 2295 27583 2301
rect 27525 2292 27537 2295
rect 26568 2264 27537 2292
rect 26568 2252 26574 2264
rect 27525 2261 27537 2264
rect 27571 2261 27583 2295
rect 27525 2255 27583 2261
rect 28537 2295 28595 2301
rect 28537 2261 28549 2295
rect 28583 2261 28595 2295
rect 28537 2255 28595 2261
rect 28994 2252 29000 2304
rect 29052 2292 29058 2304
rect 30009 2295 30067 2301
rect 30009 2292 30021 2295
rect 29052 2264 30021 2292
rect 29052 2252 29058 2264
rect 30009 2261 30021 2264
rect 30055 2261 30067 2295
rect 30116 2292 30144 2400
rect 30190 2388 30196 2440
rect 30248 2388 30254 2440
rect 30300 2437 30328 2468
rect 30285 2431 30343 2437
rect 30285 2397 30297 2431
rect 30331 2397 30343 2431
rect 30285 2391 30343 2397
rect 30558 2388 30564 2440
rect 30616 2428 30622 2440
rect 30653 2431 30711 2437
rect 30653 2428 30665 2431
rect 30616 2400 30665 2428
rect 30616 2388 30622 2400
rect 30653 2397 30665 2400
rect 30699 2397 30711 2431
rect 30653 2391 30711 2397
rect 31018 2388 31024 2440
rect 31076 2388 31082 2440
rect 31110 2292 31116 2304
rect 30116 2264 31116 2292
rect 30009 2255 30067 2261
rect 31110 2252 31116 2264
rect 31168 2252 31174 2304
rect 31220 2301 31248 2468
rect 33134 2456 33140 2508
rect 33192 2496 33198 2508
rect 33192 2468 37504 2496
rect 33192 2456 33198 2468
rect 31386 2388 31392 2440
rect 31444 2388 31450 2440
rect 32122 2388 32128 2440
rect 32180 2388 32186 2440
rect 32214 2388 32220 2440
rect 32272 2428 32278 2440
rect 36449 2431 36507 2437
rect 36449 2428 36461 2431
rect 32272 2400 36461 2428
rect 32272 2388 32278 2400
rect 36449 2397 36461 2400
rect 36495 2397 36507 2431
rect 36449 2391 36507 2397
rect 36814 2388 36820 2440
rect 36872 2388 36878 2440
rect 37476 2437 37504 2468
rect 37844 2437 37872 2536
rect 38378 2524 38384 2576
rect 38436 2524 38442 2576
rect 37461 2431 37519 2437
rect 37461 2397 37473 2431
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 37829 2431 37887 2437
rect 37829 2397 37841 2431
rect 37875 2397 37887 2431
rect 37829 2391 37887 2397
rect 38194 2388 38200 2440
rect 38252 2388 38258 2440
rect 31205 2295 31263 2301
rect 31205 2261 31217 2295
rect 31251 2261 31263 2295
rect 31205 2255 31263 2261
rect 31294 2252 31300 2304
rect 31352 2292 31358 2304
rect 32309 2295 32367 2301
rect 32309 2292 32321 2295
rect 31352 2264 32321 2292
rect 31352 2252 31358 2264
rect 32309 2261 32321 2264
rect 32355 2261 32367 2295
rect 32309 2255 32367 2261
rect 36630 2252 36636 2304
rect 36688 2252 36694 2304
rect 37001 2295 37059 2301
rect 37001 2261 37013 2295
rect 37047 2292 37059 2295
rect 37182 2292 37188 2304
rect 37047 2264 37188 2292
rect 37047 2261 37059 2264
rect 37001 2255 37059 2261
rect 37182 2252 37188 2264
rect 37240 2252 37246 2304
rect 37642 2252 37648 2304
rect 37700 2252 37706 2304
rect 38010 2252 38016 2304
rect 38068 2252 38074 2304
rect 1104 2202 38824 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 9010 2202
rect 9062 2150 9074 2202
rect 9126 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 15010 2202
rect 15062 2150 15074 2202
rect 15126 2150 15138 2202
rect 15190 2150 15202 2202
rect 15254 2150 15266 2202
rect 15318 2150 21010 2202
rect 21062 2150 21074 2202
rect 21126 2150 21138 2202
rect 21190 2150 21202 2202
rect 21254 2150 21266 2202
rect 21318 2150 27010 2202
rect 27062 2150 27074 2202
rect 27126 2150 27138 2202
rect 27190 2150 27202 2202
rect 27254 2150 27266 2202
rect 27318 2150 33010 2202
rect 33062 2150 33074 2202
rect 33126 2150 33138 2202
rect 33190 2150 33202 2202
rect 33254 2150 33266 2202
rect 33318 2150 38824 2202
rect 1104 2128 38824 2150
rect 13078 2048 13084 2100
rect 13136 2088 13142 2100
rect 24762 2088 24768 2100
rect 13136 2060 24768 2088
rect 13136 2048 13142 2060
rect 24762 2048 24768 2060
rect 24820 2048 24826 2100
rect 29546 2048 29552 2100
rect 29604 2088 29610 2100
rect 30466 2088 30472 2100
rect 29604 2060 30472 2088
rect 29604 2048 29610 2060
rect 30466 2048 30472 2060
rect 30524 2048 30530 2100
rect 32214 2088 32220 2100
rect 31726 2060 32220 2088
rect 15470 1980 15476 2032
rect 15528 2020 15534 2032
rect 15528 1992 23336 2020
rect 15528 1980 15534 1992
rect 11790 1912 11796 1964
rect 11848 1952 11854 1964
rect 22278 1952 22284 1964
rect 11848 1924 22284 1952
rect 11848 1912 11854 1924
rect 22278 1912 22284 1924
rect 22336 1912 22342 1964
rect 8478 1844 8484 1896
rect 8536 1884 8542 1896
rect 20806 1884 20812 1896
rect 8536 1856 20812 1884
rect 8536 1844 8542 1856
rect 20806 1844 20812 1856
rect 20864 1844 20870 1896
rect 23308 1884 23336 1992
rect 23382 1980 23388 2032
rect 23440 2020 23446 2032
rect 31726 2020 31754 2060
rect 32214 2048 32220 2060
rect 32272 2048 32278 2100
rect 38194 2020 38200 2032
rect 23440 1992 31754 2020
rect 35866 1992 38200 2020
rect 23440 1980 23446 1992
rect 24486 1912 24492 1964
rect 24544 1952 24550 1964
rect 35866 1952 35894 1992
rect 38194 1980 38200 1992
rect 38252 1980 38258 2032
rect 24544 1924 35894 1952
rect 24544 1912 24550 1924
rect 30282 1884 30288 1896
rect 23308 1856 30288 1884
rect 30282 1844 30288 1856
rect 30340 1844 30346 1896
rect 30466 1844 30472 1896
rect 30524 1884 30530 1896
rect 36814 1884 36820 1896
rect 30524 1856 36820 1884
rect 30524 1844 30530 1856
rect 36814 1844 36820 1856
rect 36872 1844 36878 1896
rect 13354 1776 13360 1828
rect 13412 1816 13418 1828
rect 24394 1816 24400 1828
rect 13412 1788 24400 1816
rect 13412 1776 13418 1788
rect 24394 1776 24400 1788
rect 24452 1776 24458 1828
rect 28626 1776 28632 1828
rect 28684 1816 28690 1828
rect 32122 1816 32128 1828
rect 28684 1788 32128 1816
rect 28684 1776 28690 1788
rect 32122 1776 32128 1788
rect 32180 1776 32186 1828
rect 17862 1708 17868 1760
rect 17920 1748 17926 1760
rect 25958 1748 25964 1760
rect 17920 1720 25964 1748
rect 17920 1708 17926 1720
rect 25958 1708 25964 1720
rect 26016 1708 26022 1760
rect 28534 1708 28540 1760
rect 28592 1748 28598 1760
rect 35066 1748 35072 1760
rect 28592 1720 35072 1748
rect 28592 1708 28598 1720
rect 35066 1708 35072 1720
rect 35124 1708 35130 1760
rect 14458 1640 14464 1692
rect 14516 1680 14522 1692
rect 23658 1680 23664 1692
rect 14516 1652 23664 1680
rect 14516 1640 14522 1652
rect 23658 1640 23664 1652
rect 23716 1640 23722 1692
rect 20346 1572 20352 1624
rect 20404 1612 20410 1624
rect 27706 1612 27712 1624
rect 20404 1584 27712 1612
rect 20404 1572 20410 1584
rect 27706 1572 27712 1584
rect 27764 1572 27770 1624
rect 22830 1504 22836 1556
rect 22888 1544 22894 1556
rect 30466 1544 30472 1556
rect 22888 1516 30472 1544
rect 22888 1504 22894 1516
rect 30466 1504 30472 1516
rect 30524 1504 30530 1556
rect 22370 1368 22376 1420
rect 22428 1408 22434 1420
rect 23014 1408 23020 1420
rect 22428 1380 23020 1408
rect 22428 1368 22434 1380
rect 23014 1368 23020 1380
rect 23072 1368 23078 1420
rect 11514 1300 11520 1352
rect 11572 1340 11578 1352
rect 18046 1340 18052 1352
rect 11572 1312 18052 1340
rect 11572 1300 11578 1312
rect 18046 1300 18052 1312
rect 18104 1300 18110 1352
rect 29638 1300 29644 1352
rect 29696 1340 29702 1352
rect 34790 1340 34796 1352
rect 29696 1312 34796 1340
rect 29696 1300 29702 1312
rect 34790 1300 34796 1312
rect 34848 1300 34854 1352
rect 26602 1232 26608 1284
rect 26660 1272 26666 1284
rect 33686 1272 33692 1284
rect 26660 1244 33692 1272
rect 26660 1232 26666 1244
rect 33686 1232 33692 1244
rect 33744 1232 33750 1284
rect 16022 484 16028 536
rect 16080 524 16086 536
rect 25314 524 25320 536
rect 16080 496 25320 524
rect 16080 484 16086 496
rect 25314 484 25320 496
rect 25372 484 25378 536
rect 25590 416 25596 468
rect 25648 456 25654 468
rect 33502 456 33508 468
rect 25648 428 33508 456
rect 25648 416 25654 428
rect 33502 416 33508 428
rect 33560 416 33566 468
rect 21450 348 21456 400
rect 21508 388 21514 400
rect 32306 388 32312 400
rect 21508 360 32312 388
rect 21508 348 21514 360
rect 32306 348 32312 360
rect 32364 348 32370 400
rect 16574 280 16580 332
rect 16632 320 16638 332
rect 27798 320 27804 332
rect 16632 292 27804 320
rect 16632 280 16638 292
rect 27798 280 27804 292
rect 27856 280 27862 332
rect 12986 212 12992 264
rect 13044 252 13050 264
rect 26418 252 26424 264
rect 13044 224 26424 252
rect 13044 212 13050 224
rect 26418 212 26424 224
rect 26476 212 26482 264
rect 13814 144 13820 196
rect 13872 184 13878 196
rect 28350 184 28356 196
rect 13872 156 28356 184
rect 13872 144 13878 156
rect 28350 144 28356 156
rect 28408 144 28414 196
rect 14182 76 14188 128
rect 14240 116 14246 128
rect 29178 116 29184 128
rect 14240 88 29184 116
rect 14240 76 14246 88
rect 29178 76 29184 88
rect 29236 76 29242 128
rect 14458 8 14464 60
rect 14516 48 14522 60
rect 29454 48 29460 60
rect 14516 20 29460 48
rect 14516 8 14522 20
rect 29454 8 29460 20
rect 29512 8 29518 60
<< via1 >>
rect 7380 9256 7432 9308
rect 20904 9256 20956 9308
rect 20352 9188 20404 9240
rect 36176 9188 36228 9240
rect 14740 9120 14792 9172
rect 23388 9120 23440 9172
rect 12900 9052 12952 9104
rect 25136 9052 25188 9104
rect 17224 8984 17276 9036
rect 23664 8984 23716 9036
rect 18512 8916 18564 8968
rect 37832 8916 37884 8968
rect 5540 8848 5592 8900
rect 16764 8848 16816 8900
rect 16948 8848 17000 8900
rect 25872 8848 25924 8900
rect 10784 8780 10836 8832
rect 16488 8780 16540 8832
rect 18420 8780 18472 8832
rect 26516 8780 26568 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 9010 8678 9062 8730
rect 9074 8678 9126 8730
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 15010 8678 15062 8730
rect 15074 8678 15126 8730
rect 15138 8678 15190 8730
rect 15202 8678 15254 8730
rect 15266 8678 15318 8730
rect 21010 8678 21062 8730
rect 21074 8678 21126 8730
rect 21138 8678 21190 8730
rect 21202 8678 21254 8730
rect 21266 8678 21318 8730
rect 27010 8678 27062 8730
rect 27074 8678 27126 8730
rect 27138 8678 27190 8730
rect 27202 8678 27254 8730
rect 27266 8678 27318 8730
rect 33010 8678 33062 8730
rect 33074 8678 33126 8730
rect 33138 8678 33190 8730
rect 33202 8678 33254 8730
rect 33266 8678 33318 8730
rect 1492 8576 1544 8628
rect 3424 8576 3476 8628
rect 5172 8576 5224 8628
rect 7012 8576 7064 8628
rect 8852 8576 8904 8628
rect 10692 8576 10744 8628
rect 12532 8576 12584 8628
rect 14372 8576 14424 8628
rect 16212 8576 16264 8628
rect 18052 8576 18104 8628
rect 19892 8576 19944 8628
rect 5540 8483 5592 8492
rect 5540 8449 5549 8483
rect 5549 8449 5583 8483
rect 5583 8449 5592 8483
rect 5540 8440 5592 8449
rect 7380 8483 7432 8492
rect 7380 8449 7389 8483
rect 7389 8449 7423 8483
rect 7423 8449 7432 8483
rect 7380 8440 7432 8449
rect 10784 8440 10836 8492
rect 17224 8508 17276 8560
rect 17316 8508 17368 8560
rect 21640 8576 21692 8628
rect 21732 8576 21784 8628
rect 23572 8576 23624 8628
rect 25412 8576 25464 8628
rect 27344 8576 27396 8628
rect 29092 8576 29144 8628
rect 30932 8576 30984 8628
rect 32772 8576 32824 8628
rect 34612 8576 34664 8628
rect 36360 8619 36412 8628
rect 36360 8585 36369 8619
rect 36369 8585 36403 8619
rect 36403 8585 36412 8619
rect 36360 8576 36412 8585
rect 36452 8576 36504 8628
rect 12900 8483 12952 8492
rect 12900 8449 12909 8483
rect 12909 8449 12943 8483
rect 12943 8449 12952 8483
rect 12900 8440 12952 8449
rect 14740 8483 14792 8492
rect 14740 8449 14749 8483
rect 14749 8449 14783 8483
rect 14783 8449 14792 8483
rect 14740 8440 14792 8449
rect 16948 8483 17000 8492
rect 16948 8449 16957 8483
rect 16957 8449 16991 8483
rect 16991 8449 17000 8483
rect 16948 8440 17000 8449
rect 18420 8483 18472 8492
rect 18420 8449 18429 8483
rect 18429 8449 18463 8483
rect 18463 8449 18472 8483
rect 18420 8440 18472 8449
rect 25688 8508 25740 8560
rect 38292 8576 38344 8628
rect 38936 8508 38988 8560
rect 22100 8483 22152 8492
rect 22100 8449 22109 8483
rect 22109 8449 22143 8483
rect 22143 8449 22152 8483
rect 22100 8440 22152 8449
rect 22376 8372 22428 8424
rect 25780 8483 25832 8492
rect 25780 8449 25789 8483
rect 25789 8449 25823 8483
rect 25823 8449 25832 8483
rect 25780 8440 25832 8449
rect 27620 8483 27672 8492
rect 27620 8449 27629 8483
rect 27629 8449 27663 8483
rect 27663 8449 27672 8483
rect 27620 8440 27672 8449
rect 30748 8440 30800 8492
rect 31300 8483 31352 8492
rect 31300 8449 31309 8483
rect 31309 8449 31343 8483
rect 31343 8449 31352 8483
rect 31300 8440 31352 8449
rect 34244 8440 34296 8492
rect 34980 8483 35032 8492
rect 34980 8449 34989 8483
rect 34989 8449 35023 8483
rect 35023 8449 35032 8483
rect 34980 8440 35032 8449
rect 36176 8483 36228 8492
rect 36176 8449 36185 8483
rect 36185 8449 36219 8483
rect 36219 8449 36228 8483
rect 36176 8440 36228 8449
rect 36820 8483 36872 8492
rect 36820 8449 36829 8483
rect 36829 8449 36863 8483
rect 36863 8449 36872 8483
rect 36820 8440 36872 8449
rect 28816 8372 28868 8424
rect 17316 8304 17368 8356
rect 19708 8304 19760 8356
rect 37832 8483 37884 8492
rect 37832 8449 37841 8483
rect 37841 8449 37875 8483
rect 37875 8449 37884 8483
rect 37832 8440 37884 8449
rect 37556 8372 37608 8424
rect 38752 8304 38804 8356
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 13950 8134 14002 8186
rect 14014 8134 14066 8186
rect 14078 8134 14130 8186
rect 14142 8134 14194 8186
rect 14206 8134 14258 8186
rect 19950 8134 20002 8186
rect 20014 8134 20066 8186
rect 20078 8134 20130 8186
rect 20142 8134 20194 8186
rect 20206 8134 20258 8186
rect 25950 8134 26002 8186
rect 26014 8134 26066 8186
rect 26078 8134 26130 8186
rect 26142 8134 26194 8186
rect 26206 8134 26258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 37950 8134 38002 8186
rect 38014 8134 38066 8186
rect 38078 8134 38130 8186
rect 38142 8134 38194 8186
rect 38206 8134 38258 8186
rect 36912 8075 36964 8084
rect 36912 8041 36921 8075
rect 36921 8041 36955 8075
rect 36955 8041 36964 8075
rect 36912 8032 36964 8041
rect 37280 8075 37332 8084
rect 37280 8041 37289 8075
rect 37289 8041 37323 8075
rect 37323 8041 37332 8075
rect 37280 8032 37332 8041
rect 37648 8075 37700 8084
rect 37648 8041 37657 8075
rect 37657 8041 37691 8075
rect 37691 8041 37700 8075
rect 37648 8032 37700 8041
rect 25228 7964 25280 8016
rect 26884 7964 26936 8016
rect 16856 7896 16908 7948
rect 15660 7828 15712 7880
rect 17684 7760 17736 7812
rect 18696 7760 18748 7812
rect 18788 7760 18840 7812
rect 37096 7871 37148 7880
rect 37096 7837 37105 7871
rect 37105 7837 37139 7871
rect 37139 7837 37148 7871
rect 37096 7828 37148 7837
rect 37464 7871 37516 7880
rect 37464 7837 37473 7871
rect 37473 7837 37507 7871
rect 37507 7837 37516 7871
rect 37464 7828 37516 7837
rect 18236 7692 18288 7744
rect 19248 7692 19300 7744
rect 20536 7692 20588 7744
rect 25228 7692 25280 7744
rect 38016 7735 38068 7744
rect 38016 7701 38025 7735
rect 38025 7701 38059 7735
rect 38059 7701 38068 7735
rect 38016 7692 38068 7701
rect 38384 7735 38436 7744
rect 38384 7701 38393 7735
rect 38393 7701 38427 7735
rect 38427 7701 38436 7735
rect 38384 7692 38436 7701
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 9010 7590 9062 7642
rect 9074 7590 9126 7642
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 15010 7590 15062 7642
rect 15074 7590 15126 7642
rect 15138 7590 15190 7642
rect 15202 7590 15254 7642
rect 15266 7590 15318 7642
rect 21010 7590 21062 7642
rect 21074 7590 21126 7642
rect 21138 7590 21190 7642
rect 21202 7590 21254 7642
rect 21266 7590 21318 7642
rect 27010 7590 27062 7642
rect 27074 7590 27126 7642
rect 27138 7590 27190 7642
rect 27202 7590 27254 7642
rect 27266 7590 27318 7642
rect 33010 7590 33062 7642
rect 33074 7590 33126 7642
rect 33138 7590 33190 7642
rect 33202 7590 33254 7642
rect 33266 7590 33318 7642
rect 14924 7488 14976 7540
rect 16856 7531 16908 7540
rect 16856 7497 16865 7531
rect 16865 7497 16899 7531
rect 16899 7497 16908 7531
rect 16856 7488 16908 7497
rect 17040 7531 17092 7540
rect 17040 7497 17049 7531
rect 17049 7497 17083 7531
rect 17083 7497 17092 7531
rect 17040 7488 17092 7497
rect 14832 7420 14884 7472
rect 15292 7395 15344 7404
rect 15292 7361 15301 7395
rect 15301 7361 15335 7395
rect 15335 7361 15344 7395
rect 17684 7531 17736 7540
rect 17684 7497 17693 7531
rect 17693 7497 17727 7531
rect 17727 7497 17736 7531
rect 17684 7488 17736 7497
rect 18052 7531 18104 7540
rect 18052 7497 18061 7531
rect 18061 7497 18095 7531
rect 18095 7497 18104 7531
rect 18052 7488 18104 7497
rect 18696 7420 18748 7472
rect 15292 7352 15344 7361
rect 14648 7284 14700 7336
rect 15660 7259 15712 7268
rect 15660 7225 15669 7259
rect 15669 7225 15703 7259
rect 15703 7225 15712 7259
rect 15660 7216 15712 7225
rect 16488 7216 16540 7268
rect 18236 7395 18288 7404
rect 18236 7361 18245 7395
rect 18245 7361 18279 7395
rect 18279 7361 18288 7395
rect 18236 7352 18288 7361
rect 18328 7216 18380 7268
rect 18512 7352 18564 7404
rect 18604 7395 18656 7404
rect 18604 7361 18613 7395
rect 18613 7361 18647 7395
rect 18647 7361 18656 7395
rect 18604 7352 18656 7361
rect 19248 7395 19300 7404
rect 19248 7361 19257 7395
rect 19257 7361 19291 7395
rect 19291 7361 19300 7395
rect 19248 7352 19300 7361
rect 19524 7395 19576 7404
rect 19524 7361 19533 7395
rect 19533 7361 19567 7395
rect 19567 7361 19576 7395
rect 19524 7352 19576 7361
rect 19800 7395 19852 7404
rect 19800 7361 19809 7395
rect 19809 7361 19843 7395
rect 19843 7361 19852 7395
rect 19800 7352 19852 7361
rect 20536 7395 20588 7404
rect 20536 7361 20545 7395
rect 20545 7361 20579 7395
rect 20579 7361 20588 7395
rect 20536 7352 20588 7361
rect 21364 7352 21416 7404
rect 18512 7216 18564 7268
rect 18788 7259 18840 7268
rect 18788 7225 18797 7259
rect 18797 7225 18831 7259
rect 18831 7225 18840 7259
rect 18788 7216 18840 7225
rect 15936 7191 15988 7200
rect 15936 7157 15945 7191
rect 15945 7157 15979 7191
rect 15979 7157 15988 7191
rect 15936 7148 15988 7157
rect 16764 7148 16816 7200
rect 19708 7259 19760 7268
rect 19708 7225 19717 7259
rect 19717 7225 19751 7259
rect 19751 7225 19760 7259
rect 19708 7216 19760 7225
rect 21456 7216 21508 7268
rect 21824 7531 21876 7540
rect 21824 7497 21833 7531
rect 21833 7497 21867 7531
rect 21867 7497 21876 7531
rect 21824 7488 21876 7497
rect 22376 7531 22428 7540
rect 22376 7497 22385 7531
rect 22385 7497 22419 7531
rect 22419 7497 22428 7531
rect 22376 7488 22428 7497
rect 32588 7488 32640 7540
rect 38476 7488 38528 7540
rect 23388 7420 23440 7472
rect 25320 7420 25372 7472
rect 21824 7352 21876 7404
rect 22284 7352 22336 7404
rect 22560 7395 22612 7404
rect 22560 7361 22569 7395
rect 22569 7361 22603 7395
rect 22603 7361 22612 7395
rect 22560 7352 22612 7361
rect 24124 7352 24176 7404
rect 26148 7420 26200 7472
rect 26424 7420 26476 7472
rect 25596 7352 25648 7404
rect 26148 7284 26200 7336
rect 33968 7352 34020 7404
rect 26608 7284 26660 7336
rect 26884 7284 26936 7336
rect 31852 7284 31904 7336
rect 37280 7284 37332 7336
rect 37464 7216 37516 7268
rect 20076 7148 20128 7200
rect 20260 7148 20312 7200
rect 20904 7148 20956 7200
rect 23664 7191 23716 7200
rect 23664 7157 23673 7191
rect 23673 7157 23707 7191
rect 23707 7157 23716 7191
rect 23664 7148 23716 7157
rect 25136 7148 25188 7200
rect 25320 7148 25372 7200
rect 25872 7148 25924 7200
rect 26516 7148 26568 7200
rect 38384 7191 38436 7200
rect 38384 7157 38393 7191
rect 38393 7157 38427 7191
rect 38427 7157 38436 7191
rect 38384 7148 38436 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 13950 7046 14002 7098
rect 14014 7046 14066 7098
rect 14078 7046 14130 7098
rect 14142 7046 14194 7098
rect 14206 7046 14258 7098
rect 19950 7046 20002 7098
rect 20014 7046 20066 7098
rect 20078 7046 20130 7098
rect 20142 7046 20194 7098
rect 20206 7046 20258 7098
rect 25950 7046 26002 7098
rect 26014 7046 26066 7098
rect 26078 7046 26130 7098
rect 26142 7046 26194 7098
rect 26206 7046 26258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 37950 7046 38002 7098
rect 38014 7046 38066 7098
rect 38078 7046 38130 7098
rect 38142 7046 38194 7098
rect 38206 7046 38258 7098
rect 15936 6944 15988 6996
rect 37096 6944 37148 6996
rect 1308 6808 1360 6860
rect 7840 6808 7892 6860
rect 7748 6740 7800 6792
rect 7472 6672 7524 6724
rect 8392 6783 8444 6792
rect 8392 6749 8401 6783
rect 8401 6749 8435 6783
rect 8435 6749 8444 6783
rect 8392 6740 8444 6749
rect 8208 6672 8260 6724
rect 7564 6647 7616 6656
rect 7564 6613 7573 6647
rect 7573 6613 7607 6647
rect 7607 6613 7616 6647
rect 7564 6604 7616 6613
rect 7656 6604 7708 6656
rect 8484 6604 8536 6656
rect 8576 6647 8628 6656
rect 8576 6613 8585 6647
rect 8585 6613 8619 6647
rect 8619 6613 8628 6647
rect 8576 6604 8628 6613
rect 8668 6604 8720 6656
rect 9496 6740 9548 6792
rect 10324 6783 10376 6792
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 10324 6740 10376 6749
rect 9404 6604 9456 6656
rect 9956 6604 10008 6656
rect 11796 6672 11848 6724
rect 15752 6851 15804 6860
rect 15752 6817 15761 6851
rect 15761 6817 15795 6851
rect 15795 6817 15804 6851
rect 15752 6808 15804 6817
rect 34152 6740 34204 6792
rect 20076 6672 20128 6724
rect 38200 6783 38252 6792
rect 38200 6749 38209 6783
rect 38209 6749 38243 6783
rect 38243 6749 38252 6783
rect 38200 6740 38252 6749
rect 11612 6604 11664 6656
rect 16120 6647 16172 6656
rect 16120 6613 16129 6647
rect 16129 6613 16163 6647
rect 16163 6613 16172 6647
rect 16120 6604 16172 6613
rect 20168 6647 20220 6656
rect 20168 6613 20177 6647
rect 20177 6613 20211 6647
rect 20211 6613 20220 6647
rect 20168 6604 20220 6613
rect 25688 6604 25740 6656
rect 38016 6647 38068 6656
rect 38016 6613 38025 6647
rect 38025 6613 38059 6647
rect 38059 6613 38068 6647
rect 38016 6604 38068 6613
rect 38384 6647 38436 6656
rect 38384 6613 38393 6647
rect 38393 6613 38427 6647
rect 38427 6613 38436 6647
rect 38384 6604 38436 6613
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 9010 6502 9062 6554
rect 9074 6502 9126 6554
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 15010 6502 15062 6554
rect 15074 6502 15126 6554
rect 15138 6502 15190 6554
rect 15202 6502 15254 6554
rect 15266 6502 15318 6554
rect 21010 6502 21062 6554
rect 21074 6502 21126 6554
rect 21138 6502 21190 6554
rect 21202 6502 21254 6554
rect 21266 6502 21318 6554
rect 27010 6502 27062 6554
rect 27074 6502 27126 6554
rect 27138 6502 27190 6554
rect 27202 6502 27254 6554
rect 27266 6502 27318 6554
rect 33010 6502 33062 6554
rect 33074 6502 33126 6554
rect 33138 6502 33190 6554
rect 33202 6502 33254 6554
rect 33266 6502 33318 6554
rect 6920 6400 6972 6452
rect 8668 6400 8720 6452
rect 10968 6400 11020 6452
rect 7564 6332 7616 6384
rect 11060 6332 11112 6384
rect 16672 6443 16724 6452
rect 16672 6409 16681 6443
rect 16681 6409 16715 6443
rect 16715 6409 16724 6443
rect 16672 6400 16724 6409
rect 20076 6400 20128 6452
rect 20168 6400 20220 6452
rect 37280 6400 37332 6452
rect 38384 6443 38436 6452
rect 38384 6409 38393 6443
rect 38393 6409 38427 6443
rect 38427 6409 38436 6443
rect 38384 6400 38436 6409
rect 15200 6332 15252 6384
rect 19064 6332 19116 6384
rect 6644 6264 6696 6316
rect 9496 6264 9548 6316
rect 9588 6307 9640 6316
rect 9588 6273 9597 6307
rect 9597 6273 9631 6307
rect 9631 6273 9640 6307
rect 9588 6264 9640 6273
rect 8300 6196 8352 6248
rect 10508 6264 10560 6316
rect 11336 6264 11388 6316
rect 16580 6264 16632 6316
rect 17776 6264 17828 6316
rect 11244 6196 11296 6248
rect 18788 6196 18840 6248
rect 6092 6128 6144 6180
rect 10508 6128 10560 6180
rect 10600 6171 10652 6180
rect 10600 6137 10609 6171
rect 10609 6137 10643 6171
rect 10643 6137 10652 6171
rect 10600 6128 10652 6137
rect 11152 6128 11204 6180
rect 18880 6128 18932 6180
rect 20352 6128 20404 6180
rect 37832 6128 37884 6180
rect 7196 6060 7248 6112
rect 8208 6060 8260 6112
rect 8576 6060 8628 6112
rect 12624 6060 12676 6112
rect 12716 6060 12768 6112
rect 19708 6060 19760 6112
rect 39120 6060 39172 6112
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 13950 5958 14002 6010
rect 14014 5958 14066 6010
rect 14078 5958 14130 6010
rect 14142 5958 14194 6010
rect 14206 5958 14258 6010
rect 19950 5958 20002 6010
rect 20014 5958 20066 6010
rect 20078 5958 20130 6010
rect 20142 5958 20194 6010
rect 20206 5958 20258 6010
rect 25950 5958 26002 6010
rect 26014 5958 26066 6010
rect 26078 5958 26130 6010
rect 26142 5958 26194 6010
rect 26206 5958 26258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 37950 5958 38002 6010
rect 38014 5958 38066 6010
rect 38078 5958 38130 6010
rect 38142 5958 38194 6010
rect 38206 5958 38258 6010
rect 7656 5856 7708 5908
rect 11152 5856 11204 5908
rect 6368 5788 6420 5840
rect 10324 5788 10376 5840
rect 10600 5788 10652 5840
rect 18512 5856 18564 5908
rect 18696 5899 18748 5908
rect 18696 5865 18705 5899
rect 18705 5865 18739 5899
rect 18739 5865 18748 5899
rect 18696 5856 18748 5865
rect 19064 5899 19116 5908
rect 19064 5865 19073 5899
rect 19073 5865 19107 5899
rect 19107 5865 19116 5899
rect 19064 5856 19116 5865
rect 22100 5856 22152 5908
rect 34244 5899 34296 5908
rect 34244 5865 34253 5899
rect 34253 5865 34287 5899
rect 34287 5865 34296 5899
rect 34244 5856 34296 5865
rect 34980 5856 35032 5908
rect 36820 5856 36872 5908
rect 37556 5856 37608 5908
rect 4160 5720 4212 5772
rect 9588 5720 9640 5772
rect 11060 5720 11112 5772
rect 14280 5831 14332 5840
rect 14280 5797 14289 5831
rect 14289 5797 14323 5831
rect 14323 5797 14332 5831
rect 14280 5788 14332 5797
rect 15200 5788 15252 5840
rect 22928 5788 22980 5840
rect 4988 5652 5040 5704
rect 4712 5584 4764 5636
rect 11428 5652 11480 5704
rect 19340 5720 19392 5772
rect 21364 5720 21416 5772
rect 13176 5695 13228 5704
rect 13176 5661 13185 5695
rect 13185 5661 13219 5695
rect 13219 5661 13228 5695
rect 13176 5652 13228 5661
rect 13544 5695 13596 5704
rect 13544 5661 13553 5695
rect 13553 5661 13587 5695
rect 13587 5661 13596 5695
rect 13544 5652 13596 5661
rect 13636 5652 13688 5704
rect 34520 5788 34572 5840
rect 38384 5831 38436 5840
rect 38384 5797 38393 5831
rect 38393 5797 38427 5831
rect 38427 5797 38436 5831
rect 38384 5788 38436 5797
rect 36176 5720 36228 5772
rect 36452 5652 36504 5704
rect 36728 5652 36780 5704
rect 37004 5695 37056 5704
rect 37004 5661 37013 5695
rect 37013 5661 37047 5695
rect 37047 5661 37056 5695
rect 37004 5652 37056 5661
rect 37832 5695 37884 5704
rect 37832 5661 37841 5695
rect 37841 5661 37875 5695
rect 37875 5661 37884 5695
rect 37832 5652 37884 5661
rect 11244 5584 11296 5636
rect 12716 5584 12768 5636
rect 16580 5584 16632 5636
rect 20444 5584 20496 5636
rect 13084 5559 13136 5568
rect 13084 5525 13093 5559
rect 13093 5525 13127 5559
rect 13127 5525 13136 5559
rect 13084 5516 13136 5525
rect 13360 5559 13412 5568
rect 13360 5525 13369 5559
rect 13369 5525 13403 5559
rect 13403 5525 13412 5559
rect 13360 5516 13412 5525
rect 21548 5516 21600 5568
rect 38016 5559 38068 5568
rect 38016 5525 38025 5559
rect 38025 5525 38059 5559
rect 38059 5525 38068 5559
rect 38016 5516 38068 5525
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 9010 5414 9062 5466
rect 9074 5414 9126 5466
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 15010 5414 15062 5466
rect 15074 5414 15126 5466
rect 15138 5414 15190 5466
rect 15202 5414 15254 5466
rect 15266 5414 15318 5466
rect 21010 5414 21062 5466
rect 21074 5414 21126 5466
rect 21138 5414 21190 5466
rect 21202 5414 21254 5466
rect 21266 5414 21318 5466
rect 27010 5414 27062 5466
rect 27074 5414 27126 5466
rect 27138 5414 27190 5466
rect 27202 5414 27254 5466
rect 27266 5414 27318 5466
rect 33010 5414 33062 5466
rect 33074 5414 33126 5466
rect 33138 5414 33190 5466
rect 33202 5414 33254 5466
rect 33266 5414 33318 5466
rect 4436 5312 4488 5364
rect 17316 5312 17368 5364
rect 17408 5355 17460 5364
rect 17408 5321 17417 5355
rect 17417 5321 17451 5355
rect 17451 5321 17460 5355
rect 17408 5312 17460 5321
rect 17776 5355 17828 5364
rect 17776 5321 17785 5355
rect 17785 5321 17819 5355
rect 17819 5321 17828 5355
rect 17776 5312 17828 5321
rect 20352 5312 20404 5364
rect 31116 5312 31168 5364
rect 31300 5312 31352 5364
rect 38384 5355 38436 5364
rect 38384 5321 38393 5355
rect 38393 5321 38427 5355
rect 38427 5321 38436 5355
rect 38384 5312 38436 5321
rect 11152 5244 11204 5296
rect 12440 5244 12492 5296
rect 5264 5176 5316 5228
rect 5356 5176 5408 5228
rect 10508 5176 10560 5228
rect 20536 5244 20588 5296
rect 5816 5108 5868 5160
rect 12164 5108 12216 5160
rect 5540 5040 5592 5092
rect 4620 5015 4672 5024
rect 4620 4981 4629 5015
rect 4629 4981 4663 5015
rect 4663 4981 4672 5015
rect 4620 4972 4672 4981
rect 7564 5040 7616 5092
rect 10232 5040 10284 5092
rect 17776 5176 17828 5228
rect 35992 5176 36044 5228
rect 24860 5108 24912 5160
rect 27896 5108 27948 5160
rect 31392 5108 31444 5160
rect 19616 5040 19668 5092
rect 5724 5015 5776 5024
rect 5724 4981 5733 5015
rect 5733 4981 5767 5015
rect 5767 4981 5776 5015
rect 5724 4972 5776 4981
rect 13820 4972 13872 5024
rect 14372 4972 14424 5024
rect 17592 4972 17644 5024
rect 22836 5015 22888 5024
rect 22836 4981 22845 5015
rect 22845 4981 22879 5015
rect 22879 4981 22888 5015
rect 22836 4972 22888 4981
rect 23204 5015 23256 5024
rect 23204 4981 23213 5015
rect 23213 4981 23247 5015
rect 23247 4981 23256 5015
rect 23204 4972 23256 4981
rect 23296 5015 23348 5024
rect 23296 4981 23305 5015
rect 23305 4981 23339 5015
rect 23339 4981 23348 5015
rect 23296 4972 23348 4981
rect 28172 4972 28224 5024
rect 30564 4972 30616 5024
rect 39120 4972 39172 5024
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 13950 4870 14002 4922
rect 14014 4870 14066 4922
rect 14078 4870 14130 4922
rect 14142 4870 14194 4922
rect 14206 4870 14258 4922
rect 19950 4870 20002 4922
rect 20014 4870 20066 4922
rect 20078 4870 20130 4922
rect 20142 4870 20194 4922
rect 20206 4870 20258 4922
rect 25950 4870 26002 4922
rect 26014 4870 26066 4922
rect 26078 4870 26130 4922
rect 26142 4870 26194 4922
rect 26206 4870 26258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 37950 4870 38002 4922
rect 38014 4870 38066 4922
rect 38078 4870 38130 4922
rect 38142 4870 38194 4922
rect 38206 4870 38258 4922
rect 4436 4811 4488 4820
rect 4436 4777 4445 4811
rect 4445 4777 4479 4811
rect 4479 4777 4488 4811
rect 4436 4768 4488 4777
rect 4620 4768 4672 4820
rect 11520 4768 11572 4820
rect 15476 4811 15528 4820
rect 15476 4777 15485 4811
rect 15485 4777 15519 4811
rect 15519 4777 15528 4811
rect 15476 4768 15528 4777
rect 17868 4768 17920 4820
rect 19616 4811 19668 4820
rect 19616 4777 19625 4811
rect 19625 4777 19659 4811
rect 19659 4777 19668 4811
rect 19616 4768 19668 4777
rect 2780 4700 2832 4752
rect 5356 4700 5408 4752
rect 11060 4700 11112 4752
rect 21640 4700 21692 4752
rect 27528 4768 27580 4820
rect 27620 4768 27672 4820
rect 30748 4811 30800 4820
rect 30748 4777 30757 4811
rect 30757 4777 30791 4811
rect 30791 4777 30800 4811
rect 30748 4768 30800 4777
rect 30840 4768 30892 4820
rect 35348 4768 35400 4820
rect 13820 4632 13872 4684
rect 25504 4700 25556 4752
rect 26332 4700 26384 4752
rect 31116 4700 31168 4752
rect 38200 4700 38252 4752
rect 38384 4743 38436 4752
rect 38384 4709 38393 4743
rect 38393 4709 38427 4743
rect 38427 4709 38436 4743
rect 38384 4700 38436 4709
rect 2872 4564 2924 4616
rect 9680 4564 9732 4616
rect 15568 4564 15620 4616
rect 23204 4632 23256 4684
rect 21364 4607 21416 4616
rect 21364 4573 21373 4607
rect 21373 4573 21407 4607
rect 21407 4573 21416 4607
rect 21364 4564 21416 4573
rect 5724 4496 5776 4548
rect 13820 4496 13872 4548
rect 15476 4496 15528 4548
rect 17868 4428 17920 4480
rect 21640 4496 21692 4548
rect 25688 4564 25740 4616
rect 23756 4471 23808 4480
rect 23756 4437 23765 4471
rect 23765 4437 23799 4471
rect 23799 4437 23808 4471
rect 23756 4428 23808 4437
rect 24216 4428 24268 4480
rect 29000 4607 29052 4616
rect 29000 4573 29009 4607
rect 29009 4573 29043 4607
rect 29043 4573 29052 4607
rect 29000 4564 29052 4573
rect 27804 4496 27856 4548
rect 30840 4564 30892 4616
rect 35624 4632 35676 4684
rect 27896 4471 27948 4480
rect 27896 4437 27905 4471
rect 27905 4437 27939 4471
rect 27939 4437 27948 4471
rect 27896 4428 27948 4437
rect 28172 4471 28224 4480
rect 28172 4437 28181 4471
rect 28181 4437 28215 4471
rect 28215 4437 28224 4471
rect 28172 4428 28224 4437
rect 28816 4471 28868 4480
rect 28816 4437 28825 4471
rect 28825 4437 28859 4471
rect 28859 4437 28868 4471
rect 28816 4428 28868 4437
rect 38016 4471 38068 4480
rect 38016 4437 38025 4471
rect 38025 4437 38059 4471
rect 38059 4437 38068 4471
rect 38016 4428 38068 4437
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 9010 4326 9062 4378
rect 9074 4326 9126 4378
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 15010 4326 15062 4378
rect 15074 4326 15126 4378
rect 15138 4326 15190 4378
rect 15202 4326 15254 4378
rect 15266 4326 15318 4378
rect 21010 4326 21062 4378
rect 21074 4326 21126 4378
rect 21138 4326 21190 4378
rect 21202 4326 21254 4378
rect 21266 4326 21318 4378
rect 27010 4326 27062 4378
rect 27074 4326 27126 4378
rect 27138 4326 27190 4378
rect 27202 4326 27254 4378
rect 27266 4326 27318 4378
rect 33010 4326 33062 4378
rect 33074 4326 33126 4378
rect 33138 4326 33190 4378
rect 33202 4326 33254 4378
rect 33266 4326 33318 4378
rect 572 4224 624 4276
rect 19432 4224 19484 4276
rect 19616 4224 19668 4276
rect 5724 4156 5776 4208
rect 15844 4156 15896 4208
rect 19800 4156 19852 4208
rect 22376 4156 22428 4208
rect 23756 4224 23808 4276
rect 24400 4156 24452 4208
rect 29000 4156 29052 4208
rect 29644 4156 29696 4208
rect 3608 4088 3660 4140
rect 9404 4088 9456 4140
rect 20720 4088 20772 4140
rect 7656 4020 7708 4072
rect 19340 4020 19392 4072
rect 23848 4020 23900 4072
rect 24952 4020 25004 4072
rect 27804 4088 27856 4140
rect 28356 4131 28408 4140
rect 28356 4097 28365 4131
rect 28365 4097 28399 4131
rect 28399 4097 28408 4131
rect 28356 4088 28408 4097
rect 29184 4131 29236 4140
rect 29184 4097 29193 4131
rect 29193 4097 29227 4131
rect 29227 4097 29236 4131
rect 29184 4088 29236 4097
rect 28540 4020 28592 4072
rect 29552 4020 29604 4072
rect 30288 4020 30340 4072
rect 38200 4131 38252 4140
rect 38200 4097 38209 4131
rect 38209 4097 38243 4131
rect 38243 4097 38252 4131
rect 38200 4088 38252 4097
rect 31300 4020 31352 4072
rect 37464 4020 37516 4072
rect 3056 3927 3108 3936
rect 3056 3893 3065 3927
rect 3065 3893 3099 3927
rect 3099 3893 3108 3927
rect 3056 3884 3108 3893
rect 5632 3884 5684 3936
rect 19340 3884 19392 3936
rect 20536 3884 20588 3936
rect 22008 3995 22060 4004
rect 22008 3961 22017 3995
rect 22017 3961 22051 3995
rect 22051 3961 22060 3995
rect 22008 3952 22060 3961
rect 23480 3952 23532 4004
rect 25412 3952 25464 4004
rect 25780 3952 25832 4004
rect 28264 3952 28316 4004
rect 30472 3952 30524 4004
rect 38384 3995 38436 4004
rect 38384 3961 38393 3995
rect 38393 3961 38427 3995
rect 38427 3961 38436 3995
rect 38384 3952 38436 3961
rect 23204 3884 23256 3936
rect 25044 3884 25096 3936
rect 25872 3927 25924 3936
rect 25872 3893 25881 3927
rect 25881 3893 25915 3927
rect 25915 3893 25924 3927
rect 25872 3884 25924 3893
rect 26424 3927 26476 3936
rect 26424 3893 26433 3927
rect 26433 3893 26467 3927
rect 26467 3893 26476 3927
rect 26424 3884 26476 3893
rect 26700 3927 26752 3936
rect 26700 3893 26709 3927
rect 26709 3893 26743 3927
rect 26743 3893 26752 3927
rect 26700 3884 26752 3893
rect 27436 3884 27488 3936
rect 27896 3927 27948 3936
rect 27896 3893 27905 3927
rect 27905 3893 27939 3927
rect 27939 3893 27948 3927
rect 27896 3884 27948 3893
rect 28632 3884 28684 3936
rect 28816 3884 28868 3936
rect 29460 3884 29512 3936
rect 30012 3927 30064 3936
rect 30012 3893 30021 3927
rect 30021 3893 30055 3927
rect 30055 3893 30064 3927
rect 30012 3884 30064 3893
rect 30196 3884 30248 3936
rect 30380 3884 30432 3936
rect 30840 3927 30892 3936
rect 30840 3893 30849 3927
rect 30849 3893 30883 3927
rect 30883 3893 30892 3927
rect 30840 3884 30892 3893
rect 31116 3884 31168 3936
rect 39120 3884 39172 3936
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 13950 3782 14002 3834
rect 14014 3782 14066 3834
rect 14078 3782 14130 3834
rect 14142 3782 14194 3834
rect 14206 3782 14258 3834
rect 19950 3782 20002 3834
rect 20014 3782 20066 3834
rect 20078 3782 20130 3834
rect 20142 3782 20194 3834
rect 20206 3782 20258 3834
rect 25950 3782 26002 3834
rect 26014 3782 26066 3834
rect 26078 3782 26130 3834
rect 26142 3782 26194 3834
rect 26206 3782 26258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 37950 3782 38002 3834
rect 38014 3782 38066 3834
rect 38078 3782 38130 3834
rect 38142 3782 38194 3834
rect 38206 3782 38258 3834
rect 23480 3680 23532 3732
rect 23664 3680 23716 3732
rect 25872 3680 25924 3732
rect 28632 3680 28684 3732
rect 28724 3680 28776 3732
rect 31024 3680 31076 3732
rect 3056 3612 3108 3664
rect 15384 3612 15436 3664
rect 20352 3612 20404 3664
rect 20720 3612 20772 3664
rect 21732 3612 21784 3664
rect 21824 3655 21876 3664
rect 21824 3621 21833 3655
rect 21833 3621 21867 3655
rect 21867 3621 21876 3655
rect 21824 3612 21876 3621
rect 23480 3544 23532 3596
rect 3424 3476 3476 3528
rect 8852 3476 8904 3528
rect 16856 3519 16908 3528
rect 16856 3485 16865 3519
rect 16865 3485 16899 3519
rect 16899 3485 16908 3519
rect 16856 3476 16908 3485
rect 16948 3476 17000 3528
rect 17776 3519 17828 3528
rect 17776 3485 17785 3519
rect 17785 3485 17819 3519
rect 17819 3485 17828 3519
rect 17776 3476 17828 3485
rect 19340 3476 19392 3528
rect 20720 3476 20772 3528
rect 21640 3519 21692 3528
rect 21640 3485 21649 3519
rect 21649 3485 21683 3519
rect 21683 3485 21692 3519
rect 21640 3476 21692 3485
rect 21732 3476 21784 3528
rect 23664 3519 23716 3528
rect 23664 3485 23673 3519
rect 23673 3485 23707 3519
rect 23707 3485 23716 3519
rect 23664 3476 23716 3485
rect 9588 3408 9640 3460
rect 24400 3519 24452 3528
rect 24400 3485 24409 3519
rect 24409 3485 24443 3519
rect 24443 3485 24452 3519
rect 24400 3476 24452 3485
rect 29276 3519 29328 3528
rect 29276 3485 29285 3519
rect 29285 3485 29319 3519
rect 29319 3485 29328 3519
rect 29276 3476 29328 3485
rect 3976 3383 4028 3392
rect 3976 3349 3985 3383
rect 3985 3349 4019 3383
rect 4019 3349 4028 3383
rect 3976 3340 4028 3349
rect 12624 3340 12676 3392
rect 17684 3340 17736 3392
rect 17960 3383 18012 3392
rect 17960 3349 17969 3383
rect 17969 3349 18003 3383
rect 18003 3349 18012 3383
rect 17960 3340 18012 3349
rect 20628 3340 20680 3392
rect 21732 3340 21784 3392
rect 22744 3340 22796 3392
rect 22836 3383 22888 3392
rect 22836 3349 22845 3383
rect 22845 3349 22879 3383
rect 22879 3349 22888 3383
rect 22836 3340 22888 3349
rect 23020 3383 23072 3392
rect 23020 3349 23029 3383
rect 23029 3349 23063 3383
rect 23063 3349 23072 3383
rect 23020 3340 23072 3349
rect 23112 3340 23164 3392
rect 29644 3408 29696 3460
rect 38384 3655 38436 3664
rect 38384 3621 38393 3655
rect 38393 3621 38427 3655
rect 38427 3621 38436 3655
rect 38384 3612 38436 3621
rect 35900 3544 35952 3596
rect 37924 3408 37976 3460
rect 24492 3340 24544 3392
rect 25320 3340 25372 3392
rect 28908 3383 28960 3392
rect 28908 3349 28917 3383
rect 28917 3349 28951 3383
rect 28951 3349 28960 3383
rect 28908 3340 28960 3349
rect 29552 3383 29604 3392
rect 29552 3349 29561 3383
rect 29561 3349 29595 3383
rect 29595 3349 29604 3383
rect 29552 3340 29604 3349
rect 29828 3383 29880 3392
rect 29828 3349 29837 3383
rect 29837 3349 29871 3383
rect 29871 3349 29880 3383
rect 29828 3340 29880 3349
rect 30288 3340 30340 3392
rect 38016 3383 38068 3392
rect 38016 3349 38025 3383
rect 38025 3349 38059 3383
rect 38059 3349 38068 3383
rect 38016 3340 38068 3349
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 9010 3238 9062 3290
rect 9074 3238 9126 3290
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 15010 3238 15062 3290
rect 15074 3238 15126 3290
rect 15138 3238 15190 3290
rect 15202 3238 15254 3290
rect 15266 3238 15318 3290
rect 21010 3238 21062 3290
rect 21074 3238 21126 3290
rect 21138 3238 21190 3290
rect 21202 3238 21254 3290
rect 21266 3238 21318 3290
rect 27010 3238 27062 3290
rect 27074 3238 27126 3290
rect 27138 3238 27190 3290
rect 27202 3238 27254 3290
rect 27266 3238 27318 3290
rect 33010 3238 33062 3290
rect 33074 3238 33126 3290
rect 33138 3238 33190 3290
rect 33202 3238 33254 3290
rect 33266 3238 33318 3290
rect 10968 3136 11020 3188
rect 21640 3136 21692 3188
rect 23296 3136 23348 3188
rect 8300 3068 8352 3120
rect 16948 3068 17000 3120
rect 8576 3000 8628 3052
rect 17776 3068 17828 3120
rect 17960 3068 18012 3120
rect 27068 3136 27120 3188
rect 23480 3068 23532 3120
rect 10784 2932 10836 2984
rect 13636 2932 13688 2984
rect 3976 2864 4028 2916
rect 18604 3043 18656 3052
rect 18604 3009 18613 3043
rect 18613 3009 18647 3043
rect 18647 3009 18656 3043
rect 18604 3000 18656 3009
rect 19708 3000 19760 3052
rect 17684 2932 17736 2984
rect 19248 2932 19300 2984
rect 17592 2864 17644 2916
rect 21548 2932 21600 2984
rect 22376 3043 22428 3052
rect 22376 3009 22385 3043
rect 22385 3009 22419 3043
rect 22419 3009 22428 3043
rect 22376 3000 22428 3009
rect 23848 3043 23900 3052
rect 23848 3009 23857 3043
rect 23857 3009 23891 3043
rect 23891 3009 23900 3043
rect 23848 3000 23900 3009
rect 24860 3000 24912 3052
rect 23204 2932 23256 2984
rect 27436 3043 27488 3052
rect 27436 3009 27445 3043
rect 27445 3009 27479 3043
rect 27479 3009 27488 3043
rect 27436 3000 27488 3009
rect 29552 3136 29604 3188
rect 29644 3136 29696 3188
rect 29828 3068 29880 3120
rect 30380 3000 30432 3052
rect 30564 3000 30616 3052
rect 22836 2864 22888 2916
rect 25872 2864 25924 2916
rect 26700 2932 26752 2984
rect 37464 3043 37516 3052
rect 37464 3009 37473 3043
rect 37473 3009 37507 3043
rect 37507 3009 37516 3043
rect 37464 3000 37516 3009
rect 38384 3179 38436 3188
rect 38384 3145 38393 3179
rect 38393 3145 38427 3179
rect 38427 3145 38436 3179
rect 38384 3136 38436 3145
rect 37924 3000 37976 3052
rect 31300 2864 31352 2916
rect 11244 2796 11296 2848
rect 11612 2796 11664 2848
rect 17408 2796 17460 2848
rect 18512 2796 18564 2848
rect 19340 2796 19392 2848
rect 22652 2796 22704 2848
rect 23204 2796 23256 2848
rect 23756 2796 23808 2848
rect 24860 2796 24912 2848
rect 25688 2796 25740 2848
rect 26884 2796 26936 2848
rect 28172 2796 28224 2848
rect 28448 2796 28500 2848
rect 29276 2796 29328 2848
rect 30380 2796 30432 2848
rect 30932 2796 30984 2848
rect 37832 2796 37884 2848
rect 39120 2796 39172 2848
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 13950 2694 14002 2746
rect 14014 2694 14066 2746
rect 14078 2694 14130 2746
rect 14142 2694 14194 2746
rect 14206 2694 14258 2746
rect 19950 2694 20002 2746
rect 20014 2694 20066 2746
rect 20078 2694 20130 2746
rect 20142 2694 20194 2746
rect 20206 2694 20258 2746
rect 25950 2694 26002 2746
rect 26014 2694 26066 2746
rect 26078 2694 26130 2746
rect 26142 2694 26194 2746
rect 26206 2694 26258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 37950 2694 38002 2746
rect 38014 2694 38066 2746
rect 38078 2694 38130 2746
rect 38142 2694 38194 2746
rect 38206 2694 38258 2746
rect 14280 2592 14332 2644
rect 7564 2524 7616 2576
rect 9496 2456 9548 2508
rect 15384 2388 15436 2440
rect 17316 2431 17368 2440
rect 17316 2397 17325 2431
rect 17325 2397 17359 2431
rect 17359 2397 17368 2431
rect 17316 2388 17368 2397
rect 13820 2320 13872 2372
rect 18052 2431 18104 2440
rect 18052 2397 18061 2431
rect 18061 2397 18095 2431
rect 18095 2397 18104 2431
rect 18052 2388 18104 2397
rect 18880 2524 18932 2576
rect 19616 2524 19668 2576
rect 18604 2456 18656 2508
rect 21824 2592 21876 2644
rect 22468 2592 22520 2644
rect 21548 2524 21600 2576
rect 18788 2431 18840 2440
rect 18788 2397 18797 2431
rect 18797 2397 18831 2431
rect 18831 2397 18840 2431
rect 18788 2388 18840 2397
rect 19248 2431 19300 2440
rect 19248 2397 19257 2431
rect 19257 2397 19291 2431
rect 19291 2397 19300 2431
rect 19248 2388 19300 2397
rect 19616 2431 19668 2440
rect 19616 2397 19625 2431
rect 19625 2397 19659 2431
rect 19659 2397 19668 2431
rect 19616 2388 19668 2397
rect 20444 2388 20496 2440
rect 20536 2388 20588 2440
rect 20812 2388 20864 2440
rect 22192 2431 22244 2440
rect 22192 2397 22201 2431
rect 22201 2397 22235 2431
rect 22235 2397 22244 2431
rect 22192 2388 22244 2397
rect 22284 2388 22336 2440
rect 22100 2320 22152 2372
rect 23480 2592 23532 2644
rect 24676 2592 24728 2644
rect 26148 2592 26200 2644
rect 26332 2592 26384 2644
rect 26792 2592 26844 2644
rect 27988 2592 28040 2644
rect 29828 2592 29880 2644
rect 24032 2524 24084 2576
rect 25136 2524 25188 2576
rect 26240 2524 26292 2576
rect 27344 2524 27396 2576
rect 28724 2524 28776 2576
rect 30104 2524 30156 2576
rect 22928 2431 22980 2440
rect 22928 2397 22937 2431
rect 22937 2397 22971 2431
rect 22971 2397 22980 2431
rect 22928 2388 22980 2397
rect 23020 2388 23072 2440
rect 23664 2431 23716 2440
rect 23664 2397 23673 2431
rect 23673 2397 23707 2431
rect 23707 2397 23716 2431
rect 23664 2388 23716 2397
rect 24400 2431 24452 2440
rect 24400 2397 24409 2431
rect 24409 2397 24443 2431
rect 24443 2397 24452 2431
rect 24400 2388 24452 2397
rect 24768 2431 24820 2440
rect 24768 2397 24777 2431
rect 24777 2397 24811 2431
rect 24811 2397 24820 2431
rect 24768 2388 24820 2397
rect 25412 2456 25464 2508
rect 25504 2431 25556 2440
rect 25504 2397 25513 2431
rect 25513 2397 25547 2431
rect 25547 2397 25556 2431
rect 25504 2388 25556 2397
rect 25780 2388 25832 2440
rect 25964 2388 26016 2440
rect 30012 2456 30064 2508
rect 30472 2567 30524 2576
rect 30472 2533 30481 2567
rect 30481 2533 30515 2567
rect 30515 2533 30524 2567
rect 30472 2524 30524 2533
rect 30656 2524 30708 2576
rect 33508 2524 33560 2576
rect 27068 2388 27120 2440
rect 27712 2431 27764 2440
rect 27712 2397 27721 2431
rect 27721 2397 27755 2431
rect 27755 2397 27764 2431
rect 27712 2388 27764 2397
rect 27896 2388 27948 2440
rect 28816 2388 28868 2440
rect 28908 2388 28960 2440
rect 17132 2295 17184 2304
rect 17132 2261 17141 2295
rect 17141 2261 17175 2295
rect 17175 2261 17184 2295
rect 17132 2252 17184 2261
rect 17684 2252 17736 2304
rect 17960 2252 18012 2304
rect 18236 2295 18288 2304
rect 18236 2261 18245 2295
rect 18245 2261 18279 2295
rect 18279 2261 18288 2295
rect 18236 2252 18288 2261
rect 18788 2252 18840 2304
rect 19064 2252 19116 2304
rect 19616 2252 19668 2304
rect 19892 2252 19944 2304
rect 20168 2295 20220 2304
rect 20168 2261 20177 2295
rect 20177 2261 20211 2295
rect 20211 2261 20220 2295
rect 20168 2252 20220 2261
rect 20444 2252 20496 2304
rect 20720 2252 20772 2304
rect 20996 2252 21048 2304
rect 21364 2252 21416 2304
rect 22468 2252 22520 2304
rect 22928 2252 22980 2304
rect 23020 2252 23072 2304
rect 24308 2320 24360 2372
rect 25412 2320 25464 2372
rect 27620 2320 27672 2372
rect 26516 2252 26568 2304
rect 29000 2252 29052 2304
rect 30196 2431 30248 2440
rect 30196 2397 30205 2431
rect 30205 2397 30239 2431
rect 30239 2397 30248 2431
rect 30196 2388 30248 2397
rect 30564 2388 30616 2440
rect 31024 2431 31076 2440
rect 31024 2397 31033 2431
rect 31033 2397 31067 2431
rect 31067 2397 31076 2431
rect 31024 2388 31076 2397
rect 31116 2252 31168 2304
rect 33140 2456 33192 2508
rect 31392 2431 31444 2440
rect 31392 2397 31401 2431
rect 31401 2397 31435 2431
rect 31435 2397 31444 2431
rect 31392 2388 31444 2397
rect 32128 2431 32180 2440
rect 32128 2397 32137 2431
rect 32137 2397 32171 2431
rect 32171 2397 32180 2431
rect 32128 2388 32180 2397
rect 32220 2388 32272 2440
rect 36820 2431 36872 2440
rect 36820 2397 36829 2431
rect 36829 2397 36863 2431
rect 36863 2397 36872 2431
rect 36820 2388 36872 2397
rect 38384 2567 38436 2576
rect 38384 2533 38393 2567
rect 38393 2533 38427 2567
rect 38427 2533 38436 2567
rect 38384 2524 38436 2533
rect 38200 2431 38252 2440
rect 38200 2397 38209 2431
rect 38209 2397 38243 2431
rect 38243 2397 38252 2431
rect 38200 2388 38252 2397
rect 31300 2252 31352 2304
rect 36636 2295 36688 2304
rect 36636 2261 36645 2295
rect 36645 2261 36679 2295
rect 36679 2261 36688 2295
rect 36636 2252 36688 2261
rect 37188 2252 37240 2304
rect 37648 2295 37700 2304
rect 37648 2261 37657 2295
rect 37657 2261 37691 2295
rect 37691 2261 37700 2295
rect 37648 2252 37700 2261
rect 38016 2295 38068 2304
rect 38016 2261 38025 2295
rect 38025 2261 38059 2295
rect 38059 2261 38068 2295
rect 38016 2252 38068 2261
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 9010 2150 9062 2202
rect 9074 2150 9126 2202
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 15010 2150 15062 2202
rect 15074 2150 15126 2202
rect 15138 2150 15190 2202
rect 15202 2150 15254 2202
rect 15266 2150 15318 2202
rect 21010 2150 21062 2202
rect 21074 2150 21126 2202
rect 21138 2150 21190 2202
rect 21202 2150 21254 2202
rect 21266 2150 21318 2202
rect 27010 2150 27062 2202
rect 27074 2150 27126 2202
rect 27138 2150 27190 2202
rect 27202 2150 27254 2202
rect 27266 2150 27318 2202
rect 33010 2150 33062 2202
rect 33074 2150 33126 2202
rect 33138 2150 33190 2202
rect 33202 2150 33254 2202
rect 33266 2150 33318 2202
rect 13084 2048 13136 2100
rect 24768 2048 24820 2100
rect 29552 2048 29604 2100
rect 30472 2048 30524 2100
rect 15476 1980 15528 2032
rect 11796 1912 11848 1964
rect 22284 1912 22336 1964
rect 8484 1844 8536 1896
rect 20812 1844 20864 1896
rect 23388 1980 23440 2032
rect 32220 2048 32272 2100
rect 24492 1912 24544 1964
rect 38200 1980 38252 2032
rect 30288 1844 30340 1896
rect 30472 1844 30524 1896
rect 36820 1844 36872 1896
rect 13360 1776 13412 1828
rect 24400 1776 24452 1828
rect 28632 1776 28684 1828
rect 32128 1776 32180 1828
rect 17868 1708 17920 1760
rect 25964 1708 26016 1760
rect 28540 1708 28592 1760
rect 35072 1708 35124 1760
rect 14464 1640 14516 1692
rect 23664 1640 23716 1692
rect 20352 1572 20404 1624
rect 27712 1572 27764 1624
rect 22836 1504 22888 1556
rect 30472 1504 30524 1556
rect 22376 1368 22428 1420
rect 23020 1368 23072 1420
rect 11520 1300 11572 1352
rect 18052 1300 18104 1352
rect 29644 1300 29696 1352
rect 34796 1300 34848 1352
rect 26608 1232 26660 1284
rect 33692 1232 33744 1284
rect 16028 484 16080 536
rect 25320 484 25372 536
rect 25596 416 25648 468
rect 33508 416 33560 468
rect 21456 348 21508 400
rect 32312 348 32364 400
rect 16580 280 16632 332
rect 27804 280 27856 332
rect 12992 212 13044 264
rect 26424 212 26476 264
rect 13820 144 13872 196
rect 28356 144 28408 196
rect 14188 76 14240 128
rect 29184 76 29236 128
rect 14464 8 14516 60
rect 29460 8 29512 60
<< metal2 >>
rect 1490 11096 1546 11152
rect 3330 11096 3386 11152
rect 5170 11096 5226 11152
rect 7010 11096 7066 11152
rect 8850 11096 8906 11152
rect 10690 11096 10746 11152
rect 12530 11096 12586 11152
rect 14370 11096 14426 11152
rect 16210 11096 16266 11152
rect 18050 11096 18106 11152
rect 19890 11096 19946 11152
rect 21730 11096 21786 11152
rect 23570 11096 23626 11152
rect 25410 11096 25466 11152
rect 27250 11096 27306 11152
rect 29090 11096 29146 11152
rect 30930 11096 30986 11152
rect 32770 11096 32826 11152
rect 34610 11096 34666 11152
rect 36450 11096 36506 11152
rect 38290 11096 38346 11152
rect 1504 8634 1532 11096
rect 3344 9602 3372 11096
rect 3344 9574 3464 9602
rect 2870 8800 2926 8809
rect 2870 8735 2926 8744
rect 1492 8628 1544 8634
rect 1492 8570 1544 8576
rect 2884 8401 2912 8735
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 3436 8634 3464 9574
rect 5184 8634 5212 11096
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5552 8498 5580 8842
rect 7024 8634 7052 11096
rect 7380 9308 7432 9314
rect 7380 9250 7432 9256
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 7392 8498 7420 9250
rect 8864 8634 8892 11096
rect 9010 8732 9318 8741
rect 9010 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9176 8732
rect 9232 8730 9256 8732
rect 9312 8730 9318 8732
rect 9072 8678 9074 8730
rect 9254 8678 9256 8730
rect 9010 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9176 8678
rect 9232 8676 9256 8678
rect 9312 8676 9318 8678
rect 9010 8667 9318 8676
rect 10704 8634 10732 11096
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10796 8498 10824 8774
rect 12544 8634 12572 11096
rect 12900 9104 12952 9110
rect 12900 9046 12952 9052
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12912 8498 12940 9046
rect 14384 8634 14412 11096
rect 14646 9344 14702 9353
rect 14646 9279 14702 9288
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 2870 8392 2926 8401
rect 2870 8327 2926 8336
rect 1766 8256 1822 8265
rect 1766 8191 1822 8200
rect 1780 7313 1808 8191
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 13950 8188 14258 8197
rect 13950 8186 13956 8188
rect 14012 8186 14036 8188
rect 14092 8186 14116 8188
rect 14172 8186 14196 8188
rect 14252 8186 14258 8188
rect 14012 8134 14014 8186
rect 14194 8134 14196 8186
rect 13950 8132 13956 8134
rect 14012 8132 14036 8134
rect 14092 8132 14116 8134
rect 14172 8132 14196 8134
rect 14252 8132 14258 8134
rect 13950 8123 14258 8132
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 9010 7644 9318 7653
rect 9010 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9176 7644
rect 9232 7642 9256 7644
rect 9312 7642 9318 7644
rect 9072 7590 9074 7642
rect 9254 7590 9256 7642
rect 9010 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9176 7590
rect 9232 7588 9256 7590
rect 9312 7588 9318 7590
rect 9010 7579 9318 7588
rect 14660 7342 14688 9279
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 14752 8498 14780 9114
rect 14830 9072 14886 9081
rect 14830 9007 14886 9016
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14844 7478 14872 9007
rect 15010 8732 15318 8741
rect 15010 8730 15016 8732
rect 15072 8730 15096 8732
rect 15152 8730 15176 8732
rect 15232 8730 15256 8732
rect 15312 8730 15318 8732
rect 15072 8678 15074 8730
rect 15254 8678 15256 8730
rect 15010 8676 15016 8678
rect 15072 8676 15096 8678
rect 15152 8676 15176 8678
rect 15232 8676 15256 8678
rect 15312 8676 15318 8678
rect 15010 8667 15318 8676
rect 16224 8634 16252 11096
rect 17224 9036 17276 9042
rect 17224 8978 17276 8984
rect 16764 8900 16816 8906
rect 16764 8842 16816 8848
rect 16948 8900 17000 8906
rect 16948 8842 17000 8848
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 14922 8392 14978 8401
rect 14922 8327 14978 8336
rect 14936 7546 14964 8327
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 15010 7644 15318 7653
rect 15010 7642 15016 7644
rect 15072 7642 15096 7644
rect 15152 7642 15176 7644
rect 15232 7642 15256 7644
rect 15312 7642 15318 7644
rect 15072 7590 15074 7642
rect 15254 7590 15256 7642
rect 15010 7588 15016 7590
rect 15072 7588 15096 7590
rect 15152 7588 15176 7590
rect 15232 7588 15256 7590
rect 15312 7588 15318 7590
rect 15010 7579 15318 7588
rect 14924 7540 14976 7546
rect 14924 7482 14976 7488
rect 14832 7472 14884 7478
rect 14832 7414 14884 7420
rect 15290 7440 15346 7449
rect 15290 7375 15292 7384
rect 15344 7375 15346 7384
rect 15292 7346 15344 7352
rect 14648 7336 14700 7342
rect 1766 7304 1822 7313
rect 14648 7278 14700 7284
rect 15672 7274 15700 7822
rect 16500 7274 16528 8774
rect 1766 7239 1822 7248
rect 15660 7268 15712 7274
rect 15660 7210 15712 7216
rect 16488 7268 16540 7274
rect 16488 7210 16540 7216
rect 16776 7206 16804 8842
rect 16960 8498 16988 8842
rect 17236 8566 17264 8978
rect 18064 8634 18092 11096
rect 19798 9616 19854 9625
rect 19798 9551 19854 9560
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18420 8832 18472 8838
rect 18420 8774 18472 8780
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 17224 8560 17276 8566
rect 17038 8528 17094 8537
rect 16948 8492 17000 8498
rect 17224 8502 17276 8508
rect 17316 8560 17368 8566
rect 17316 8502 17368 8508
rect 17038 8463 17094 8472
rect 16948 8434 17000 8440
rect 16856 7948 16908 7954
rect 16856 7890 16908 7896
rect 16868 7546 16896 7890
rect 17052 7546 17080 8463
rect 17328 8362 17356 8502
rect 18432 8498 18460 8774
rect 18420 8492 18472 8498
rect 18420 8434 18472 8440
rect 17316 8356 17368 8362
rect 17316 8298 17368 8304
rect 18234 7984 18290 7993
rect 18234 7919 18290 7928
rect 18050 7848 18106 7857
rect 17684 7812 17736 7818
rect 18050 7783 18106 7792
rect 17684 7754 17736 7760
rect 17696 7546 17724 7754
rect 18064 7546 18092 7783
rect 18248 7750 18276 7919
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 17040 7540 17092 7546
rect 17040 7482 17092 7488
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 18248 7410 18276 7686
rect 18524 7410 18552 8910
rect 19708 8356 19760 8362
rect 19708 8298 19760 8304
rect 18602 7848 18658 7857
rect 18602 7783 18658 7792
rect 18696 7812 18748 7818
rect 18616 7410 18644 7783
rect 18696 7754 18748 7760
rect 18788 7812 18840 7818
rect 18788 7754 18840 7760
rect 18708 7478 18736 7754
rect 18696 7472 18748 7478
rect 18696 7414 18748 7420
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18800 7274 18828 7754
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 19260 7410 19288 7686
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 19536 7313 19564 7346
rect 19522 7304 19578 7313
rect 18328 7268 18380 7274
rect 18512 7268 18564 7274
rect 18380 7228 18512 7256
rect 18328 7210 18380 7216
rect 18512 7210 18564 7216
rect 18788 7268 18840 7274
rect 19720 7274 19748 8298
rect 19812 7410 19840 9551
rect 19904 8634 19932 11096
rect 20904 9308 20956 9314
rect 20904 9250 20956 9256
rect 20352 9240 20404 9246
rect 20352 9182 20404 9188
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 19950 8188 20258 8197
rect 19950 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20196 8188
rect 20252 8186 20258 8188
rect 20012 8134 20014 8186
rect 20194 8134 20196 8186
rect 19950 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20196 8134
rect 20252 8132 20258 8134
rect 19950 8123 20258 8132
rect 20364 7460 20392 9182
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 20088 7432 20392 7460
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 19522 7239 19578 7248
rect 19708 7268 19760 7274
rect 18788 7210 18840 7216
rect 19708 7210 19760 7216
rect 20088 7206 20116 7432
rect 20548 7410 20576 7686
rect 20536 7404 20588 7410
rect 20536 7346 20588 7352
rect 20258 7304 20314 7313
rect 20258 7239 20314 7248
rect 20272 7206 20300 7239
rect 20916 7206 20944 9250
rect 21010 8732 21318 8741
rect 21010 8730 21016 8732
rect 21072 8730 21096 8732
rect 21152 8730 21176 8732
rect 21232 8730 21256 8732
rect 21312 8730 21318 8732
rect 21072 8678 21074 8730
rect 21254 8678 21256 8730
rect 21010 8676 21016 8678
rect 21072 8676 21096 8678
rect 21152 8676 21176 8678
rect 21232 8676 21256 8678
rect 21312 8676 21318 8678
rect 21010 8667 21318 8676
rect 21744 8634 21772 11096
rect 23388 9172 23440 9178
rect 23388 9114 23440 9120
rect 21640 8628 21692 8634
rect 21640 8570 21692 8576
rect 21732 8628 21784 8634
rect 21732 8570 21784 8576
rect 21652 7698 21680 8570
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 21652 7670 21864 7698
rect 21010 7644 21318 7653
rect 21010 7642 21016 7644
rect 21072 7642 21096 7644
rect 21152 7642 21176 7644
rect 21232 7642 21256 7644
rect 21312 7642 21318 7644
rect 21072 7590 21074 7642
rect 21254 7590 21256 7642
rect 21010 7588 21016 7590
rect 21072 7588 21096 7590
rect 21152 7588 21176 7590
rect 21232 7588 21256 7590
rect 21312 7588 21318 7590
rect 21010 7579 21318 7588
rect 21836 7546 21864 7670
rect 21824 7540 21876 7546
rect 21824 7482 21876 7488
rect 21364 7404 21416 7410
rect 21824 7404 21876 7410
rect 21416 7364 21824 7392
rect 21364 7346 21416 7352
rect 21824 7346 21876 7352
rect 21456 7268 21508 7274
rect 21456 7210 21508 7216
rect 15936 7200 15988 7206
rect 1306 7168 1362 7177
rect 15936 7142 15988 7148
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20904 7200 20956 7206
rect 20904 7142 20956 7148
rect 1306 7103 1362 7112
rect 1320 6866 1348 7103
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 13950 7100 14258 7109
rect 13950 7098 13956 7100
rect 14012 7098 14036 7100
rect 14092 7098 14116 7100
rect 14172 7098 14196 7100
rect 14252 7098 14258 7100
rect 14012 7046 14014 7098
rect 14194 7046 14196 7098
rect 13950 7044 13956 7046
rect 14012 7044 14036 7046
rect 14092 7044 14116 7046
rect 14172 7044 14196 7046
rect 14252 7044 14258 7046
rect 13950 7035 14258 7044
rect 15948 7002 15976 7142
rect 19950 7100 20258 7109
rect 19950 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20196 7100
rect 20252 7098 20258 7100
rect 20012 7046 20014 7098
rect 20194 7046 20196 7098
rect 19950 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20196 7046
rect 20252 7044 20258 7046
rect 19950 7035 20258 7044
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 15750 6896 15806 6905
rect 1308 6860 1360 6866
rect 1308 6802 1360 6808
rect 7840 6860 7892 6866
rect 15750 6831 15752 6840
rect 7840 6802 7892 6808
rect 15804 6831 15806 6840
rect 16118 6896 16174 6905
rect 16118 6831 16174 6840
rect 15752 6802 15804 6808
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7472 6724 7524 6730
rect 7472 6666 7524 6672
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6092 6180 6144 6186
rect 6092 6122 6144 6128
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 3882 5672 3938 5681
rect 3882 5607 3938 5616
rect 2870 5536 2926 5545
rect 2870 5471 2926 5480
rect 2884 5284 2912 5471
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 2884 5273 3004 5284
rect 2778 5264 2834 5273
rect 2884 5264 3018 5273
rect 2884 5256 2962 5264
rect 2778 5199 2834 5208
rect 2962 5199 3018 5208
rect 2792 5114 2820 5199
rect 2962 5128 3018 5137
rect 2792 5086 2962 5114
rect 2962 5063 3018 5072
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 2780 4752 2832 4758
rect 2780 4694 2832 4700
rect 572 4276 624 4282
rect 572 4218 624 4224
rect 584 2553 612 4218
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 570 2544 626 2553
rect 570 2479 626 2488
rect 2792 56 2820 4694
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2778 0 2834 56
rect 2884 42 2912 4558
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 3068 3670 3096 3878
rect 3056 3664 3108 3670
rect 3056 3606 3108 3612
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 3436 1714 3464 3470
rect 3344 1686 3464 1714
rect 2976 56 3096 82
rect 3344 56 3372 1686
rect 3620 56 3648 4082
rect 3896 56 3924 5607
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 3988 2922 4016 3334
rect 3976 2916 4028 2922
rect 3976 2858 4028 2864
rect 4172 56 4200 5714
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4448 4826 4476 5306
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4632 4826 4660 4966
rect 4436 4820 4488 4826
rect 4436 4762 4488 4768
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4434 4448 4490 4457
rect 4434 4383 4490 4392
rect 4448 56 4476 4383
rect 4724 56 4752 5578
rect 5000 56 5028 5646
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5276 56 5304 5170
rect 5368 4758 5396 5170
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5540 5092 5592 5098
rect 5540 5034 5592 5040
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 5552 56 5580 5034
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5736 4554 5764 4966
rect 5724 4548 5776 4554
rect 5724 4490 5776 4496
rect 5724 4208 5776 4214
rect 5724 4150 5776 4156
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5644 1465 5672 3878
rect 5736 2009 5764 4150
rect 5722 2000 5778 2009
rect 5722 1935 5778 1944
rect 5630 1456 5686 1465
rect 5630 1391 5686 1400
rect 5828 56 5856 5102
rect 6104 56 6132 6122
rect 6368 5840 6420 5846
rect 6368 5782 6420 5788
rect 6380 56 6408 5782
rect 6656 56 6684 6258
rect 6932 56 6960 6394
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 7208 56 7236 6054
rect 7484 56 7512 6666
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7576 6390 7604 6598
rect 7564 6384 7616 6390
rect 7564 6326 7616 6332
rect 7668 5914 7696 6598
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7564 5092 7616 5098
rect 7564 5034 7616 5040
rect 7576 2582 7604 5034
rect 7654 4992 7710 5001
rect 7654 4927 7710 4936
rect 7668 4078 7696 4927
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7564 2576 7616 2582
rect 7564 2518 7616 2524
rect 7760 56 7788 6734
rect 2976 54 3110 56
rect 2976 42 3004 54
rect 2884 14 3004 42
rect 3054 0 3110 54
rect 3330 0 3386 56
rect 3606 0 3662 56
rect 3882 0 3938 56
rect 4158 0 4214 56
rect 4434 0 4490 56
rect 4710 0 4766 56
rect 4986 0 5042 56
rect 5262 0 5318 56
rect 5538 0 5594 56
rect 5814 0 5870 56
rect 6090 0 6146 56
rect 6366 0 6422 56
rect 6642 0 6698 56
rect 6918 0 6974 56
rect 7194 0 7250 56
rect 7470 0 7526 56
rect 7746 0 7802 56
rect 7852 42 7880 6802
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 8220 6118 8248 6666
rect 8300 6248 8352 6254
rect 8300 6190 8352 6196
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 8312 5681 8340 6190
rect 8298 5672 8354 5681
rect 8298 5607 8354 5616
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 8404 4457 8432 6734
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 8390 4448 8446 4457
rect 8390 4383 8446 4392
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 8300 3120 8352 3126
rect 8300 3062 8352 3068
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 7944 56 8064 82
rect 8312 56 8340 3062
rect 8496 1902 8524 6598
rect 8588 6118 8616 6598
rect 8680 6458 8708 6598
rect 9010 6556 9318 6565
rect 9010 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9176 6556
rect 9232 6554 9256 6556
rect 9312 6554 9318 6556
rect 9072 6502 9074 6554
rect 9254 6502 9256 6554
rect 9010 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9176 6502
rect 9232 6500 9256 6502
rect 9312 6500 9318 6502
rect 9010 6491 9318 6500
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 9010 5468 9318 5477
rect 9010 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9176 5468
rect 9232 5466 9256 5468
rect 9312 5466 9318 5468
rect 9072 5414 9074 5466
rect 9254 5414 9256 5466
rect 9010 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9176 5414
rect 9232 5412 9256 5414
rect 9312 5412 9318 5414
rect 9010 5403 9318 5412
rect 9416 4706 9444 6598
rect 9508 6322 9536 6734
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9600 5778 9628 6258
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9968 5681 9996 6598
rect 10336 5846 10364 6734
rect 11796 6724 11848 6730
rect 11796 6666 11848 6672
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10520 6186 10548 6258
rect 10508 6180 10560 6186
rect 10508 6122 10560 6128
rect 10600 6180 10652 6186
rect 10980 6168 11008 6394
rect 11060 6384 11112 6390
rect 11112 6332 11376 6338
rect 11060 6326 11376 6332
rect 11072 6322 11376 6326
rect 11072 6316 11388 6322
rect 11072 6310 11336 6316
rect 11336 6258 11388 6264
rect 11244 6248 11296 6254
rect 11244 6190 11296 6196
rect 11152 6180 11204 6186
rect 10980 6140 11152 6168
rect 10600 6122 10652 6128
rect 11152 6122 11204 6128
rect 10612 5846 10640 6122
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 10324 5840 10376 5846
rect 10324 5782 10376 5788
rect 10600 5840 10652 5846
rect 10600 5782 10652 5788
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 9954 5672 10010 5681
rect 9954 5607 10010 5616
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10232 5092 10284 5098
rect 10232 5034 10284 5040
rect 9416 4678 9536 4706
rect 9010 4380 9318 4389
rect 9010 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9176 4380
rect 9232 4378 9256 4380
rect 9312 4378 9318 4380
rect 9072 4326 9074 4378
rect 9254 4326 9256 4378
rect 9010 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9176 4326
rect 9232 4324 9256 4326
rect 9312 4324 9318 4326
rect 9010 4315 9318 4324
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 8758 3904 8814 3913
rect 8758 3839 8814 3848
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8484 1896 8536 1902
rect 8484 1838 8536 1844
rect 8588 56 8616 2994
rect 8772 82 8800 3839
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 8864 218 8892 3470
rect 9010 3292 9318 3301
rect 9010 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9176 3292
rect 9232 3290 9256 3292
rect 9312 3290 9318 3292
rect 9072 3238 9074 3290
rect 9254 3238 9256 3290
rect 9010 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9176 3238
rect 9232 3236 9256 3238
rect 9312 3236 9318 3238
rect 9010 3227 9318 3236
rect 9010 2204 9318 2213
rect 9010 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9176 2204
rect 9232 2202 9256 2204
rect 9312 2202 9318 2204
rect 9072 2150 9074 2202
rect 9254 2150 9256 2202
rect 9010 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9176 2150
rect 9232 2148 9256 2150
rect 9312 2148 9318 2150
rect 9010 2139 9318 2148
rect 8864 190 8984 218
rect 8772 56 8892 82
rect 7944 54 8078 56
rect 7944 42 7972 54
rect 7852 14 7972 42
rect 8022 0 8078 54
rect 8298 0 8354 56
rect 8574 0 8630 56
rect 8772 54 8906 56
rect 8850 0 8906 54
rect 8956 42 8984 190
rect 9048 56 9168 82
rect 9416 56 9444 4082
rect 9508 2514 9536 4678
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9588 3460 9640 3466
rect 9588 3402 9640 3408
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9600 1737 9628 3402
rect 9586 1728 9642 1737
rect 9586 1663 9642 1672
rect 9692 56 9720 4558
rect 9954 2000 10010 2009
rect 9954 1935 10010 1944
rect 9968 56 9996 1935
rect 10244 56 10272 5034
rect 10520 56 10548 5170
rect 11072 4842 11100 5714
rect 11164 5386 11192 5850
rect 11256 5642 11284 6190
rect 11428 5704 11480 5710
rect 11428 5646 11480 5652
rect 11244 5636 11296 5642
rect 11244 5578 11296 5584
rect 11164 5358 11284 5386
rect 11152 5296 11204 5302
rect 11152 5238 11204 5244
rect 10980 4814 11100 4842
rect 10980 3890 11008 4814
rect 11060 4752 11112 4758
rect 11060 4694 11112 4700
rect 11072 4049 11100 4694
rect 11058 4040 11114 4049
rect 11058 3975 11114 3984
rect 10980 3862 11100 3890
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 10796 56 10824 2926
rect 10980 2417 11008 3130
rect 10966 2408 11022 2417
rect 10966 2343 11022 2352
rect 11072 56 11100 3862
rect 11164 3233 11192 5238
rect 11150 3224 11206 3233
rect 11150 3159 11206 3168
rect 11256 3074 11284 5358
rect 11164 3046 11284 3074
rect 11164 1601 11192 3046
rect 11244 2848 11296 2854
rect 11244 2790 11296 2796
rect 11256 2417 11284 2790
rect 11440 2774 11468 5646
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11348 2746 11468 2774
rect 11242 2408 11298 2417
rect 11242 2343 11298 2352
rect 11150 1592 11206 1601
rect 11150 1527 11206 1536
rect 11348 56 11376 2746
rect 11532 1358 11560 4762
rect 11624 2854 11652 6598
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 11610 2680 11666 2689
rect 11610 2615 11666 2624
rect 11520 1352 11572 1358
rect 11520 1294 11572 1300
rect 11624 56 11652 2615
rect 11808 1970 11836 6666
rect 16132 6662 16160 6831
rect 16670 6760 16726 6769
rect 16670 6695 16726 6704
rect 20076 6724 20128 6730
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 15010 6556 15318 6565
rect 15010 6554 15016 6556
rect 15072 6554 15096 6556
rect 15152 6554 15176 6556
rect 15232 6554 15256 6556
rect 15312 6554 15318 6556
rect 15072 6502 15074 6554
rect 15254 6502 15256 6554
rect 15010 6500 15016 6502
rect 15072 6500 15096 6502
rect 15152 6500 15176 6502
rect 15232 6500 15256 6502
rect 15312 6500 15318 6502
rect 15010 6491 15318 6500
rect 16684 6458 16712 6695
rect 20076 6666 20128 6672
rect 20088 6458 20116 6666
rect 20168 6656 20220 6662
rect 20168 6598 20220 6604
rect 20180 6458 20208 6598
rect 21010 6556 21318 6565
rect 21010 6554 21016 6556
rect 21072 6554 21096 6556
rect 21152 6554 21176 6556
rect 21232 6554 21256 6556
rect 21312 6554 21318 6556
rect 21072 6502 21074 6554
rect 21254 6502 21256 6554
rect 21010 6500 21016 6502
rect 21072 6500 21096 6502
rect 21152 6500 21176 6502
rect 21232 6500 21256 6502
rect 21312 6500 21318 6502
rect 21010 6491 21318 6500
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 20168 6452 20220 6458
rect 20168 6394 20220 6400
rect 15200 6384 15252 6390
rect 19064 6384 19116 6390
rect 15200 6326 15252 6332
rect 18694 6352 18750 6361
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12440 5296 12492 5302
rect 12440 5238 12492 5244
rect 12164 5160 12216 5166
rect 12164 5102 12216 5108
rect 11886 2544 11942 2553
rect 11886 2479 11942 2488
rect 11796 1964 11848 1970
rect 11796 1906 11848 1912
rect 11900 56 11928 2479
rect 12176 56 12204 5102
rect 12452 56 12480 5238
rect 12636 3398 12664 6054
rect 12728 5642 12756 6054
rect 13950 6012 14258 6021
rect 13950 6010 13956 6012
rect 14012 6010 14036 6012
rect 14092 6010 14116 6012
rect 14172 6010 14196 6012
rect 14252 6010 14258 6012
rect 14012 5958 14014 6010
rect 14194 5958 14196 6010
rect 13950 5956 13956 5958
rect 14012 5956 14036 5958
rect 14092 5956 14116 5958
rect 14172 5956 14196 5958
rect 14252 5956 14258 5958
rect 13950 5947 14258 5956
rect 15212 5846 15240 6326
rect 16580 6316 16632 6322
rect 16580 6258 16632 6264
rect 17776 6316 17828 6322
rect 19064 6326 19116 6332
rect 18694 6287 18750 6296
rect 17776 6258 17828 6264
rect 14280 5840 14332 5846
rect 14280 5782 14332 5788
rect 15200 5840 15252 5846
rect 15200 5782 15252 5788
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13636 5704 13688 5710
rect 13636 5646 13688 5652
rect 12716 5636 12768 5642
rect 12716 5578 12768 5584
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 13096 2106 13124 5510
rect 13188 2689 13216 5646
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 13174 2680 13230 2689
rect 13174 2615 13230 2624
rect 13084 2100 13136 2106
rect 13084 2042 13136 2048
rect 13372 1834 13400 5510
rect 13556 2553 13584 5646
rect 13648 2990 13676 5646
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13832 4690 13860 4966
rect 13950 4924 14258 4933
rect 13950 4922 13956 4924
rect 14012 4922 14036 4924
rect 14092 4922 14116 4924
rect 14172 4922 14196 4924
rect 14252 4922 14258 4924
rect 14012 4870 14014 4922
rect 14194 4870 14196 4922
rect 13950 4868 13956 4870
rect 14012 4868 14036 4870
rect 14092 4868 14116 4870
rect 14172 4868 14196 4870
rect 14252 4868 14258 4870
rect 13950 4859 14258 4868
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 13820 4548 13872 4554
rect 13820 4490 13872 4496
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 13542 2544 13598 2553
rect 13542 2479 13598 2488
rect 13832 2378 13860 4490
rect 13950 3836 14258 3845
rect 13950 3834 13956 3836
rect 14012 3834 14036 3836
rect 14092 3834 14116 3836
rect 14172 3834 14196 3836
rect 14252 3834 14258 3836
rect 14012 3782 14014 3834
rect 14194 3782 14196 3834
rect 13950 3780 13956 3782
rect 14012 3780 14036 3782
rect 14092 3780 14116 3782
rect 14172 3780 14196 3782
rect 14252 3780 14258 3782
rect 13950 3771 14258 3780
rect 13950 2748 14258 2757
rect 13950 2746 13956 2748
rect 14012 2746 14036 2748
rect 14092 2746 14116 2748
rect 14172 2746 14196 2748
rect 14252 2746 14258 2748
rect 14012 2694 14014 2746
rect 14194 2694 14196 2746
rect 13950 2692 13956 2694
rect 14012 2692 14036 2694
rect 14092 2692 14116 2694
rect 14172 2692 14196 2694
rect 14252 2692 14258 2694
rect 13950 2683 14258 2692
rect 14292 2650 14320 5782
rect 16592 5642 16620 6258
rect 17406 6216 17462 6225
rect 17406 6151 17462 6160
rect 16580 5636 16632 5642
rect 16580 5578 16632 5584
rect 15010 5468 15318 5477
rect 15010 5466 15016 5468
rect 15072 5466 15096 5468
rect 15152 5466 15176 5468
rect 15232 5466 15256 5468
rect 15312 5466 15318 5468
rect 15072 5414 15074 5466
rect 15254 5414 15256 5466
rect 15010 5412 15016 5414
rect 15072 5412 15096 5414
rect 15152 5412 15176 5414
rect 15232 5412 15256 5414
rect 15312 5412 15318 5414
rect 15010 5403 15318 5412
rect 17420 5370 17448 6151
rect 17788 5370 17816 6258
rect 18708 5914 18736 6287
rect 18788 6248 18840 6254
rect 18788 6190 18840 6196
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18696 5908 18748 5914
rect 18696 5850 18748 5856
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17408 5364 17460 5370
rect 17408 5306 17460 5312
rect 17776 5364 17828 5370
rect 17776 5306 17828 5312
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 14384 2774 14412 4966
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 15488 4554 15516 4762
rect 15568 4616 15620 4622
rect 15568 4558 15620 4564
rect 15476 4548 15528 4554
rect 15476 4490 15528 4496
rect 15010 4380 15318 4389
rect 15010 4378 15016 4380
rect 15072 4378 15096 4380
rect 15152 4378 15176 4380
rect 15232 4378 15256 4380
rect 15312 4378 15318 4380
rect 15072 4326 15074 4378
rect 15254 4326 15256 4378
rect 15010 4324 15016 4326
rect 15072 4324 15096 4326
rect 15152 4324 15176 4326
rect 15232 4324 15256 4326
rect 15312 4324 15318 4326
rect 15010 4315 15318 4324
rect 15384 3664 15436 3670
rect 15384 3606 15436 3612
rect 15010 3292 15318 3301
rect 15010 3290 15016 3292
rect 15072 3290 15096 3292
rect 15152 3290 15176 3292
rect 15232 3290 15256 3292
rect 15312 3290 15318 3292
rect 15072 3238 15074 3290
rect 15254 3238 15256 3290
rect 15010 3236 15016 3238
rect 15072 3236 15096 3238
rect 15152 3236 15176 3238
rect 15232 3236 15256 3238
rect 15312 3236 15318 3238
rect 15010 3227 15318 3236
rect 14384 2746 14504 2774
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 13360 1828 13412 1834
rect 13360 1770 13412 1776
rect 14476 1698 14504 2746
rect 15396 2446 15424 3606
rect 15384 2440 15436 2446
rect 15384 2382 15436 2388
rect 15474 2408 15530 2417
rect 15474 2343 15530 2352
rect 15010 2204 15318 2213
rect 15010 2202 15016 2204
rect 15072 2202 15096 2204
rect 15152 2202 15176 2204
rect 15232 2202 15256 2204
rect 15312 2202 15318 2204
rect 15072 2150 15074 2202
rect 15254 2150 15256 2202
rect 15010 2148 15016 2150
rect 15072 2148 15096 2150
rect 15152 2148 15176 2150
rect 15232 2148 15256 2150
rect 15312 2148 15318 2150
rect 15010 2139 15318 2148
rect 15488 2122 15516 2343
rect 15396 2094 15516 2122
rect 14464 1692 14516 1698
rect 14464 1634 14516 1640
rect 13266 640 13322 649
rect 13266 575 13322 584
rect 12714 368 12770 377
rect 12714 303 12770 312
rect 12728 56 12756 303
rect 12992 264 13044 270
rect 12992 206 13044 212
rect 13004 56 13032 206
rect 13280 56 13308 575
rect 13542 504 13598 513
rect 13542 439 13598 448
rect 13556 56 13584 439
rect 14922 232 14978 241
rect 13820 196 13872 202
rect 14922 167 14978 176
rect 13820 138 13872 144
rect 13832 56 13860 138
rect 14188 128 14240 134
rect 14108 76 14188 82
rect 14646 96 14702 105
rect 14108 70 14240 76
rect 14108 56 14228 70
rect 14384 66 14504 82
rect 14384 60 14516 66
rect 14384 56 14464 60
rect 9048 54 9182 56
rect 9048 42 9076 54
rect 8956 14 9076 42
rect 9126 0 9182 54
rect 9402 0 9458 56
rect 9678 0 9734 56
rect 9954 0 10010 56
rect 10230 0 10286 56
rect 10506 0 10562 56
rect 10782 0 10838 56
rect 11058 0 11114 56
rect 11334 0 11390 56
rect 11610 0 11666 56
rect 11886 0 11942 56
rect 12162 0 12218 56
rect 12438 0 12494 56
rect 12714 0 12770 56
rect 12990 0 13046 56
rect 13266 0 13322 56
rect 13542 0 13598 56
rect 13818 0 13874 56
rect 14094 54 14228 56
rect 14370 54 14464 56
rect 14094 0 14150 54
rect 14370 0 14426 54
rect 14464 2 14516 8
rect 14936 56 14964 167
rect 15212 56 15332 82
rect 14646 0 14702 40
rect 14922 0 14978 56
rect 15198 54 15332 56
rect 15198 0 15254 54
rect 15304 42 15332 54
rect 15396 42 15424 2094
rect 15476 2032 15528 2038
rect 15580 2009 15608 4558
rect 15842 4312 15898 4321
rect 15842 4247 15898 4256
rect 15856 4214 15884 4247
rect 15844 4208 15896 4214
rect 15844 4150 15896 4156
rect 16854 4040 16910 4049
rect 16854 3975 16910 3984
rect 16868 3534 16896 3975
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 16948 3528 17000 3534
rect 16948 3470 17000 3476
rect 15750 3360 15806 3369
rect 15750 3295 15806 3304
rect 15476 1974 15528 1980
rect 15566 2000 15622 2009
rect 15488 56 15516 1974
rect 15566 1935 15622 1944
rect 15764 56 15792 3295
rect 16960 3126 16988 3470
rect 16948 3120 17000 3126
rect 16948 3062 17000 3068
rect 17328 2446 17356 5306
rect 17774 5264 17830 5273
rect 17774 5199 17776 5208
rect 17828 5199 17830 5208
rect 17776 5170 17828 5176
rect 17866 5128 17922 5137
rect 17866 5063 17922 5072
rect 17592 5024 17644 5030
rect 17592 4966 17644 4972
rect 17604 2922 17632 4966
rect 17880 4826 17908 5063
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 17684 3392 17736 3398
rect 17684 3334 17736 3340
rect 17696 2990 17724 3334
rect 17788 3126 17816 3470
rect 17776 3120 17828 3126
rect 17776 3062 17828 3068
rect 17684 2984 17736 2990
rect 17684 2926 17736 2932
rect 17592 2916 17644 2922
rect 17592 2858 17644 2864
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 17316 2440 17368 2446
rect 17316 2382 17368 2388
rect 17132 2304 17184 2310
rect 17132 2246 17184 2252
rect 16302 1864 16358 1873
rect 16302 1799 16358 1808
rect 16028 536 16080 542
rect 16028 478 16080 484
rect 16040 56 16068 478
rect 16316 56 16344 1799
rect 16854 1728 16910 1737
rect 16854 1663 16910 1672
rect 16580 332 16632 338
rect 16580 274 16632 280
rect 16592 56 16620 274
rect 16868 56 16896 1663
rect 17144 56 17172 2246
rect 17420 56 17448 2790
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 17696 56 17724 2246
rect 17880 1766 17908 4422
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 17972 3126 18000 3334
rect 17960 3120 18012 3126
rect 17960 3062 18012 3068
rect 18524 2938 18552 5850
rect 18602 3496 18658 3505
rect 18602 3431 18658 3440
rect 18616 3058 18644 3431
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18524 2910 18644 2938
rect 18512 2848 18564 2854
rect 18512 2790 18564 2796
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 17960 2304 18012 2310
rect 17960 2246 18012 2252
rect 17868 1760 17920 1766
rect 17868 1702 17920 1708
rect 17972 56 18000 2246
rect 18064 1358 18092 2382
rect 18236 2304 18288 2310
rect 18236 2246 18288 2252
rect 18052 1352 18104 1358
rect 18052 1294 18104 1300
rect 18248 56 18276 2246
rect 18524 56 18552 2790
rect 18616 2514 18644 2910
rect 18604 2508 18656 2514
rect 18604 2450 18656 2456
rect 18800 2446 18828 6190
rect 18880 6180 18932 6186
rect 18880 6122 18932 6128
rect 18892 2582 18920 6122
rect 19076 5914 19104 6326
rect 20352 6180 20404 6186
rect 20352 6122 20404 6128
rect 19708 6112 19760 6118
rect 19708 6054 19760 6060
rect 19064 5908 19116 5914
rect 19064 5850 19116 5856
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19352 4078 19380 5714
rect 19616 5092 19668 5098
rect 19616 5034 19668 5040
rect 19628 4826 19656 5034
rect 19616 4820 19668 4826
rect 19616 4762 19668 4768
rect 19432 4276 19484 4282
rect 19432 4218 19484 4224
rect 19616 4276 19668 4282
rect 19616 4218 19668 4224
rect 19444 4162 19472 4218
rect 19628 4162 19656 4218
rect 19444 4134 19656 4162
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 19340 3936 19392 3942
rect 19340 3878 19392 3884
rect 19352 3534 19380 3878
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19720 3058 19748 6054
rect 19950 6012 20258 6021
rect 19950 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20196 6012
rect 20252 6010 20258 6012
rect 20012 5958 20014 6010
rect 20194 5958 20196 6010
rect 19950 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20196 5958
rect 20252 5956 20258 5958
rect 19950 5947 20258 5956
rect 20364 5370 20392 6122
rect 21362 5808 21418 5817
rect 21362 5743 21364 5752
rect 21416 5743 21418 5752
rect 21364 5714 21416 5720
rect 20444 5636 20496 5642
rect 20444 5578 20496 5584
rect 20352 5364 20404 5370
rect 20352 5306 20404 5312
rect 19950 4924 20258 4933
rect 19950 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20196 4924
rect 20252 4922 20258 4924
rect 20012 4870 20014 4922
rect 20194 4870 20196 4922
rect 19950 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20196 4870
rect 20252 4868 20258 4870
rect 19950 4859 20258 4868
rect 19798 4312 19854 4321
rect 19798 4247 19854 4256
rect 19812 4214 19840 4247
rect 19800 4208 19852 4214
rect 19800 4150 19852 4156
rect 19950 3836 20258 3845
rect 19950 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20196 3836
rect 20252 3834 20258 3836
rect 20012 3782 20014 3834
rect 20194 3782 20196 3834
rect 19950 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20196 3782
rect 20252 3780 20258 3782
rect 19950 3771 20258 3780
rect 20352 3664 20404 3670
rect 20352 3606 20404 3612
rect 19708 3052 19760 3058
rect 19708 2994 19760 3000
rect 19248 2984 19300 2990
rect 19248 2926 19300 2932
rect 18880 2576 18932 2582
rect 18880 2518 18932 2524
rect 19260 2446 19288 2926
rect 19340 2848 19392 2854
rect 19340 2790 19392 2796
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 19248 2440 19300 2446
rect 19248 2382 19300 2388
rect 18788 2304 18840 2310
rect 18788 2246 18840 2252
rect 19064 2304 19116 2310
rect 19064 2246 19116 2252
rect 18800 56 18828 2246
rect 19076 56 19104 2246
rect 19352 56 19380 2790
rect 19950 2748 20258 2757
rect 19950 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20196 2748
rect 20252 2746 20258 2748
rect 20012 2694 20014 2746
rect 20194 2694 20196 2746
rect 19950 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20196 2694
rect 20252 2692 20258 2694
rect 19950 2683 20258 2692
rect 19616 2576 19668 2582
rect 19616 2518 19668 2524
rect 19628 2446 19656 2518
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 19616 2304 19668 2310
rect 19616 2246 19668 2252
rect 19892 2304 19944 2310
rect 19892 2246 19944 2252
rect 20168 2304 20220 2310
rect 20168 2246 20220 2252
rect 19628 56 19656 2246
rect 19904 56 19932 2246
rect 20180 56 20208 2246
rect 20364 1630 20392 3606
rect 20456 2446 20484 5578
rect 21010 5468 21318 5477
rect 21010 5466 21016 5468
rect 21072 5466 21096 5468
rect 21152 5466 21176 5468
rect 21232 5466 21256 5468
rect 21312 5466 21318 5468
rect 21072 5414 21074 5466
rect 21254 5414 21256 5466
rect 21010 5412 21016 5414
rect 21072 5412 21096 5414
rect 21152 5412 21176 5414
rect 21232 5412 21256 5414
rect 21312 5412 21318 5414
rect 21010 5403 21318 5412
rect 20536 5296 20588 5302
rect 20536 5238 20588 5244
rect 20548 3942 20576 5238
rect 21362 4720 21418 4729
rect 21362 4655 21418 4664
rect 21376 4622 21404 4655
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 21010 4380 21318 4389
rect 21010 4378 21016 4380
rect 21072 4378 21096 4380
rect 21152 4378 21176 4380
rect 21232 4378 21256 4380
rect 21312 4378 21318 4380
rect 21072 4326 21074 4378
rect 21254 4326 21256 4378
rect 21010 4324 21016 4326
rect 21072 4324 21096 4326
rect 21152 4324 21176 4326
rect 21232 4324 21256 4326
rect 21312 4324 21318 4326
rect 21010 4315 21318 4324
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 20732 4049 20760 4082
rect 20718 4040 20774 4049
rect 20718 3975 20774 3984
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20720 3664 20772 3670
rect 20720 3606 20772 3612
rect 20732 3534 20760 3606
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 20444 2440 20496 2446
rect 20444 2382 20496 2388
rect 20536 2440 20588 2446
rect 20536 2382 20588 2388
rect 20444 2304 20496 2310
rect 20444 2246 20496 2252
rect 20352 1624 20404 1630
rect 20352 1566 20404 1572
rect 20456 56 20484 2246
rect 20548 1601 20576 2382
rect 20534 1592 20590 1601
rect 20534 1527 20590 1536
rect 20640 1193 20668 3334
rect 21010 3292 21318 3301
rect 21010 3290 21016 3292
rect 21072 3290 21096 3292
rect 21152 3290 21176 3292
rect 21232 3290 21256 3292
rect 21312 3290 21318 3292
rect 21072 3238 21074 3290
rect 21254 3238 21256 3290
rect 21010 3236 21016 3238
rect 21072 3236 21096 3238
rect 21152 3236 21176 3238
rect 21232 3236 21256 3238
rect 21312 3236 21318 3238
rect 21010 3227 21318 3236
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 20720 2304 20772 2310
rect 20720 2246 20772 2252
rect 20626 1184 20682 1193
rect 20626 1119 20682 1128
rect 20732 56 20760 2246
rect 20824 1902 20852 2382
rect 20996 2304 21048 2310
rect 20916 2264 20996 2292
rect 20812 1896 20864 1902
rect 20812 1838 20864 1844
rect 20916 1170 20944 2264
rect 20996 2246 21048 2252
rect 21364 2304 21416 2310
rect 21364 2246 21416 2252
rect 21010 2204 21318 2213
rect 21010 2202 21016 2204
rect 21072 2202 21096 2204
rect 21152 2202 21176 2204
rect 21232 2202 21256 2204
rect 21312 2202 21318 2204
rect 21072 2150 21074 2202
rect 21254 2150 21256 2202
rect 21010 2148 21016 2150
rect 21072 2148 21096 2150
rect 21152 2148 21176 2150
rect 21232 2148 21256 2150
rect 21312 2148 21318 2150
rect 21010 2139 21318 2148
rect 21376 1170 21404 2246
rect 20916 1142 21036 1170
rect 21008 56 21036 1142
rect 21284 1142 21404 1170
rect 21284 56 21312 1142
rect 21468 406 21496 7210
rect 22112 5914 22140 8434
rect 22376 8424 22428 8430
rect 22376 8366 22428 8372
rect 22388 7546 22416 8366
rect 22376 7540 22428 7546
rect 22376 7482 22428 7488
rect 23400 7478 23428 9114
rect 23584 8634 23612 11096
rect 25136 9104 25188 9110
rect 25136 9046 25188 9052
rect 23664 9036 23716 9042
rect 23664 8978 23716 8984
rect 23572 8628 23624 8634
rect 23572 8570 23624 8576
rect 23388 7472 23440 7478
rect 23388 7414 23440 7420
rect 22284 7404 22336 7410
rect 22284 7346 22336 7352
rect 22560 7404 22612 7410
rect 22560 7346 22612 7352
rect 22296 6225 22324 7346
rect 22282 6216 22338 6225
rect 22282 6151 22338 6160
rect 22100 5908 22152 5914
rect 22100 5850 22152 5856
rect 22190 5672 22246 5681
rect 22190 5607 22246 5616
rect 21548 5568 21600 5574
rect 21548 5510 21600 5516
rect 21560 2990 21588 5510
rect 21640 4752 21692 4758
rect 21640 4694 21692 4700
rect 21652 4554 21680 4694
rect 21640 4548 21692 4554
rect 21640 4490 21692 4496
rect 22006 4040 22062 4049
rect 22006 3975 22008 3984
rect 22060 3975 22062 3984
rect 22008 3946 22060 3952
rect 21732 3664 21784 3670
rect 21824 3664 21876 3670
rect 21732 3606 21784 3612
rect 21822 3632 21824 3641
rect 21876 3632 21878 3641
rect 21744 3534 21772 3606
rect 21822 3567 21878 3576
rect 21640 3528 21692 3534
rect 21640 3470 21692 3476
rect 21732 3528 21784 3534
rect 21732 3470 21784 3476
rect 21652 3194 21680 3470
rect 21732 3392 21784 3398
rect 21732 3334 21784 3340
rect 21640 3188 21692 3194
rect 21640 3130 21692 3136
rect 21548 2984 21600 2990
rect 21744 2961 21772 3334
rect 21548 2926 21600 2932
rect 21730 2952 21786 2961
rect 21730 2887 21786 2896
rect 21824 2644 21876 2650
rect 21824 2586 21876 2592
rect 21548 2576 21600 2582
rect 21548 2518 21600 2524
rect 21456 400 21508 406
rect 21456 342 21508 348
rect 21560 56 21588 2518
rect 21836 56 21864 2586
rect 22204 2446 22232 5607
rect 22376 4208 22428 4214
rect 22376 4150 22428 4156
rect 22388 3058 22416 4150
rect 22376 3052 22428 3058
rect 22376 2994 22428 3000
rect 22468 2644 22520 2650
rect 22468 2586 22520 2592
rect 22192 2440 22244 2446
rect 22192 2382 22244 2388
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 22100 2372 22152 2378
rect 22100 2314 22152 2320
rect 22112 56 22140 2314
rect 22296 1970 22324 2382
rect 22480 2310 22508 2586
rect 22468 2304 22520 2310
rect 22468 2246 22520 2252
rect 22284 1964 22336 1970
rect 22284 1906 22336 1912
rect 22572 1465 22600 7346
rect 23676 7206 23704 8978
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 23664 7200 23716 7206
rect 23664 7142 23716 7148
rect 22928 5840 22980 5846
rect 22928 5782 22980 5788
rect 22836 5024 22888 5030
rect 22836 4966 22888 4972
rect 22848 4593 22876 4966
rect 22834 4584 22890 4593
rect 22834 4519 22890 4528
rect 22744 3392 22796 3398
rect 22744 3334 22796 3340
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 22652 2848 22704 2854
rect 22652 2790 22704 2796
rect 22558 1456 22614 1465
rect 22376 1420 22428 1426
rect 22558 1391 22614 1400
rect 22376 1362 22428 1368
rect 22388 56 22416 1362
rect 22664 56 22692 2790
rect 22756 2774 22784 3334
rect 22848 2922 22876 3334
rect 22836 2916 22888 2922
rect 22836 2858 22888 2864
rect 22940 2774 22968 5782
rect 23204 5024 23256 5030
rect 23204 4966 23256 4972
rect 23296 5024 23348 5030
rect 23296 4966 23348 4972
rect 23216 4690 23244 4966
rect 23204 4684 23256 4690
rect 23204 4626 23256 4632
rect 23308 4185 23336 4966
rect 23756 4480 23808 4486
rect 23756 4422 23808 4428
rect 23768 4282 23796 4422
rect 23756 4276 23808 4282
rect 23756 4218 23808 4224
rect 23294 4176 23350 4185
rect 23294 4111 23350 4120
rect 23848 4072 23900 4078
rect 23848 4014 23900 4020
rect 23480 4004 23532 4010
rect 23480 3946 23532 3952
rect 23204 3936 23256 3942
rect 23204 3878 23256 3884
rect 23020 3392 23072 3398
rect 23020 3334 23072 3340
rect 23112 3392 23164 3398
rect 23112 3334 23164 3340
rect 23032 3097 23060 3334
rect 23018 3088 23074 3097
rect 23018 3023 23074 3032
rect 23124 2825 23152 3334
rect 23216 2990 23244 3878
rect 23492 3738 23520 3946
rect 23662 3768 23718 3777
rect 23480 3732 23532 3738
rect 23662 3703 23664 3712
rect 23480 3674 23532 3680
rect 23716 3703 23718 3712
rect 23664 3674 23716 3680
rect 23480 3596 23532 3602
rect 23480 3538 23532 3544
rect 23296 3188 23348 3194
rect 23296 3130 23348 3136
rect 23204 2984 23256 2990
rect 23204 2926 23256 2932
rect 23204 2848 23256 2854
rect 23110 2816 23166 2825
rect 22756 2746 22876 2774
rect 22940 2746 23060 2774
rect 23204 2790 23256 2796
rect 23110 2751 23166 2760
rect 22848 1562 22876 2746
rect 22926 2544 22982 2553
rect 22926 2479 22982 2488
rect 22940 2446 22968 2479
rect 23032 2446 23060 2746
rect 22928 2440 22980 2446
rect 22928 2382 22980 2388
rect 23020 2440 23072 2446
rect 23020 2382 23072 2388
rect 22928 2304 22980 2310
rect 22928 2246 22980 2252
rect 23020 2304 23072 2310
rect 23020 2246 23072 2252
rect 22836 1556 22888 1562
rect 22836 1498 22888 1504
rect 22940 56 22968 2246
rect 23032 1426 23060 2246
rect 23020 1420 23072 1426
rect 23020 1362 23072 1368
rect 23216 56 23244 2790
rect 23308 2774 23336 3130
rect 23492 3126 23520 3538
rect 23676 3534 23704 3674
rect 23664 3528 23716 3534
rect 23664 3470 23716 3476
rect 23480 3120 23532 3126
rect 23480 3062 23532 3068
rect 23860 3058 23888 4014
rect 23848 3052 23900 3058
rect 23848 2994 23900 3000
rect 23756 2848 23808 2854
rect 23756 2790 23808 2796
rect 23308 2746 23428 2774
rect 23400 2038 23428 2746
rect 23480 2644 23532 2650
rect 23480 2586 23532 2592
rect 23388 2032 23440 2038
rect 23388 1974 23440 1980
rect 23492 56 23520 2586
rect 23664 2440 23716 2446
rect 23664 2382 23716 2388
rect 23676 1698 23704 2382
rect 23664 1692 23716 1698
rect 23664 1634 23716 1640
rect 23768 56 23796 2790
rect 24032 2576 24084 2582
rect 24136 2553 24164 7346
rect 25148 7206 25176 9046
rect 25424 8634 25452 11096
rect 27264 8922 27292 11096
rect 25872 8900 25924 8906
rect 27264 8894 27384 8922
rect 25872 8842 25924 8848
rect 25412 8628 25464 8634
rect 25412 8570 25464 8576
rect 25688 8560 25740 8566
rect 25688 8502 25740 8508
rect 25228 8016 25280 8022
rect 25228 7958 25280 7964
rect 25240 7750 25268 7958
rect 25228 7744 25280 7750
rect 25228 7686 25280 7692
rect 25320 7472 25372 7478
rect 25320 7414 25372 7420
rect 25332 7206 25360 7414
rect 25596 7404 25648 7410
rect 25596 7346 25648 7352
rect 25136 7200 25188 7206
rect 25136 7142 25188 7148
rect 25320 7200 25372 7206
rect 25320 7142 25372 7148
rect 24860 5160 24912 5166
rect 24860 5102 24912 5108
rect 24216 4480 24268 4486
rect 24216 4422 24268 4428
rect 24032 2518 24084 2524
rect 24122 2544 24178 2553
rect 24044 56 24072 2518
rect 24122 2479 24178 2488
rect 24228 649 24256 4422
rect 24400 4208 24452 4214
rect 24400 4150 24452 4156
rect 24412 3534 24440 4150
rect 24400 3528 24452 3534
rect 24400 3470 24452 3476
rect 24492 3392 24544 3398
rect 24492 3334 24544 3340
rect 24400 2440 24452 2446
rect 24400 2382 24452 2388
rect 24308 2372 24360 2378
rect 24308 2314 24360 2320
rect 24214 640 24270 649
rect 24214 575 24270 584
rect 24320 56 24348 2314
rect 24412 1834 24440 2382
rect 24504 1970 24532 3334
rect 24872 3058 24900 5102
rect 25504 4752 25556 4758
rect 25504 4694 25556 4700
rect 24952 4072 25004 4078
rect 24952 4014 25004 4020
rect 24860 3052 24912 3058
rect 24860 2994 24912 3000
rect 24860 2848 24912 2854
rect 24860 2790 24912 2796
rect 24676 2644 24728 2650
rect 24596 2604 24676 2632
rect 24492 1964 24544 1970
rect 24492 1906 24544 1912
rect 24400 1828 24452 1834
rect 24400 1770 24452 1776
rect 24596 56 24624 2604
rect 24676 2586 24728 2592
rect 24768 2440 24820 2446
rect 24768 2382 24820 2388
rect 24780 2106 24808 2382
rect 24768 2100 24820 2106
rect 24768 2042 24820 2048
rect 24872 56 24900 2790
rect 24964 1737 24992 4014
rect 25412 4004 25464 4010
rect 25412 3946 25464 3952
rect 25044 3936 25096 3942
rect 25044 3878 25096 3884
rect 24950 1728 25006 1737
rect 24950 1663 25006 1672
rect 25056 377 25084 3878
rect 25320 3392 25372 3398
rect 25320 3334 25372 3340
rect 25136 2576 25188 2582
rect 25136 2518 25188 2524
rect 25042 368 25098 377
rect 25042 303 25098 312
rect 25148 56 25176 2518
rect 25332 542 25360 3334
rect 25424 2514 25452 3946
rect 25412 2508 25464 2514
rect 25412 2450 25464 2456
rect 25516 2446 25544 4694
rect 25504 2440 25556 2446
rect 25504 2382 25556 2388
rect 25412 2372 25464 2378
rect 25412 2314 25464 2320
rect 25320 536 25372 542
rect 25320 478 25372 484
rect 25424 56 25452 2314
rect 25608 474 25636 7346
rect 25700 6662 25728 8502
rect 25780 8492 25832 8498
rect 25780 8434 25832 8440
rect 25688 6656 25740 6662
rect 25688 6598 25740 6604
rect 25688 4616 25740 4622
rect 25688 4558 25740 4564
rect 25700 3890 25728 4558
rect 25792 4010 25820 8434
rect 25884 7206 25912 8842
rect 26516 8832 26568 8838
rect 26516 8774 26568 8780
rect 25950 8188 26258 8197
rect 25950 8186 25956 8188
rect 26012 8186 26036 8188
rect 26092 8186 26116 8188
rect 26172 8186 26196 8188
rect 26252 8186 26258 8188
rect 26012 8134 26014 8186
rect 26194 8134 26196 8186
rect 25950 8132 25956 8134
rect 26012 8132 26036 8134
rect 26092 8132 26116 8134
rect 26172 8132 26196 8134
rect 26252 8132 26258 8134
rect 25950 8123 26258 8132
rect 26148 7472 26200 7478
rect 26424 7472 26476 7478
rect 26238 7440 26294 7449
rect 26200 7420 26238 7426
rect 26148 7414 26238 7420
rect 26160 7398 26238 7414
rect 26424 7414 26476 7420
rect 26238 7375 26294 7384
rect 26148 7336 26200 7342
rect 26436 7290 26464 7414
rect 26200 7284 26464 7290
rect 26148 7278 26464 7284
rect 26160 7262 26464 7278
rect 26528 7206 26556 8774
rect 27010 8732 27318 8741
rect 27010 8730 27016 8732
rect 27072 8730 27096 8732
rect 27152 8730 27176 8732
rect 27232 8730 27256 8732
rect 27312 8730 27318 8732
rect 27072 8678 27074 8730
rect 27254 8678 27256 8730
rect 27010 8676 27016 8678
rect 27072 8676 27096 8678
rect 27152 8676 27176 8678
rect 27232 8676 27256 8678
rect 27312 8676 27318 8678
rect 27010 8667 27318 8676
rect 27356 8634 27384 8894
rect 29104 8634 29132 11096
rect 30944 8634 30972 11096
rect 32784 8634 32812 11096
rect 33010 8732 33318 8741
rect 33010 8730 33016 8732
rect 33072 8730 33096 8732
rect 33152 8730 33176 8732
rect 33232 8730 33256 8732
rect 33312 8730 33318 8732
rect 33072 8678 33074 8730
rect 33254 8678 33256 8730
rect 33010 8676 33016 8678
rect 33072 8676 33096 8678
rect 33152 8676 33176 8678
rect 33232 8676 33256 8678
rect 33312 8676 33318 8678
rect 33010 8667 33318 8676
rect 34624 8634 34652 11096
rect 36358 9616 36414 9625
rect 36358 9551 36414 9560
rect 36176 9240 36228 9246
rect 36176 9182 36228 9188
rect 27344 8628 27396 8634
rect 27344 8570 27396 8576
rect 29092 8628 29144 8634
rect 29092 8570 29144 8576
rect 30932 8628 30984 8634
rect 30932 8570 30984 8576
rect 32772 8628 32824 8634
rect 32772 8570 32824 8576
rect 34612 8628 34664 8634
rect 34612 8570 34664 8576
rect 36188 8498 36216 9182
rect 36372 8634 36400 9551
rect 36464 8634 36492 11096
rect 36910 9344 36966 9353
rect 36910 9279 36966 9288
rect 36360 8628 36412 8634
rect 36360 8570 36412 8576
rect 36452 8628 36504 8634
rect 36452 8570 36504 8576
rect 27620 8492 27672 8498
rect 27620 8434 27672 8440
rect 30748 8492 30800 8498
rect 30748 8434 30800 8440
rect 31300 8492 31352 8498
rect 31300 8434 31352 8440
rect 34244 8492 34296 8498
rect 34244 8434 34296 8440
rect 34980 8492 35032 8498
rect 34980 8434 35032 8440
rect 36176 8492 36228 8498
rect 36176 8434 36228 8440
rect 36820 8492 36872 8498
rect 36820 8434 36872 8440
rect 26884 8016 26936 8022
rect 26884 7958 26936 7964
rect 26896 7342 26924 7958
rect 27010 7644 27318 7653
rect 27010 7642 27016 7644
rect 27072 7642 27096 7644
rect 27152 7642 27176 7644
rect 27232 7642 27256 7644
rect 27312 7642 27318 7644
rect 27072 7590 27074 7642
rect 27254 7590 27256 7642
rect 27010 7588 27016 7590
rect 27072 7588 27096 7590
rect 27152 7588 27176 7590
rect 27232 7588 27256 7590
rect 27312 7588 27318 7590
rect 27010 7579 27318 7588
rect 26608 7336 26660 7342
rect 26608 7278 26660 7284
rect 26884 7336 26936 7342
rect 26884 7278 26936 7284
rect 25872 7200 25924 7206
rect 25872 7142 25924 7148
rect 26516 7200 26568 7206
rect 26516 7142 26568 7148
rect 25950 7100 26258 7109
rect 25950 7098 25956 7100
rect 26012 7098 26036 7100
rect 26092 7098 26116 7100
rect 26172 7098 26196 7100
rect 26252 7098 26258 7100
rect 26012 7046 26014 7098
rect 26194 7046 26196 7098
rect 25950 7044 25956 7046
rect 26012 7044 26036 7046
rect 26092 7044 26116 7046
rect 26172 7044 26196 7046
rect 26252 7044 26258 7046
rect 25950 7035 26258 7044
rect 25950 6012 26258 6021
rect 25950 6010 25956 6012
rect 26012 6010 26036 6012
rect 26092 6010 26116 6012
rect 26172 6010 26196 6012
rect 26252 6010 26258 6012
rect 26012 5958 26014 6010
rect 26194 5958 26196 6010
rect 25950 5956 25956 5958
rect 26012 5956 26036 5958
rect 26092 5956 26116 5958
rect 26172 5956 26196 5958
rect 26252 5956 26258 5958
rect 25950 5947 26258 5956
rect 25950 4924 26258 4933
rect 25950 4922 25956 4924
rect 26012 4922 26036 4924
rect 26092 4922 26116 4924
rect 26172 4922 26196 4924
rect 26252 4922 26258 4924
rect 26012 4870 26014 4922
rect 26194 4870 26196 4922
rect 25950 4868 25956 4870
rect 26012 4868 26036 4870
rect 26092 4868 26116 4870
rect 26172 4868 26196 4870
rect 26252 4868 26258 4870
rect 25950 4859 26258 4868
rect 26332 4752 26384 4758
rect 26332 4694 26384 4700
rect 25780 4004 25832 4010
rect 25780 3946 25832 3952
rect 25872 3936 25924 3942
rect 25700 3862 25820 3890
rect 25872 3878 25924 3884
rect 25688 2848 25740 2854
rect 25688 2790 25740 2796
rect 25596 468 25648 474
rect 25596 410 25648 416
rect 25700 56 25728 2790
rect 25792 2446 25820 3862
rect 25884 3738 25912 3878
rect 25950 3836 26258 3845
rect 25950 3834 25956 3836
rect 26012 3834 26036 3836
rect 26092 3834 26116 3836
rect 26172 3834 26196 3836
rect 26252 3834 26258 3836
rect 26012 3782 26014 3834
rect 26194 3782 26196 3834
rect 25950 3780 25956 3782
rect 26012 3780 26036 3782
rect 26092 3780 26116 3782
rect 26172 3780 26196 3782
rect 26252 3780 26258 3782
rect 25950 3771 26258 3780
rect 25872 3732 25924 3738
rect 25872 3674 25924 3680
rect 25872 2916 25924 2922
rect 25872 2858 25924 2864
rect 25780 2440 25832 2446
rect 25780 2382 25832 2388
rect 25884 1442 25912 2858
rect 25950 2748 26258 2757
rect 25950 2746 25956 2748
rect 26012 2746 26036 2748
rect 26092 2746 26116 2748
rect 26172 2746 26196 2748
rect 26252 2746 26258 2748
rect 26012 2694 26014 2746
rect 26194 2694 26196 2746
rect 25950 2692 25956 2694
rect 26012 2692 26036 2694
rect 26092 2692 26116 2694
rect 26172 2692 26196 2694
rect 26252 2692 26258 2694
rect 25950 2683 26258 2692
rect 26344 2650 26372 4694
rect 26424 3936 26476 3942
rect 26424 3878 26476 3884
rect 26148 2644 26200 2650
rect 26148 2586 26200 2592
rect 26332 2644 26384 2650
rect 26332 2586 26384 2592
rect 25964 2440 26016 2446
rect 25964 2382 26016 2388
rect 25976 1766 26004 2382
rect 25964 1760 26016 1766
rect 25964 1702 26016 1708
rect 25884 1414 26004 1442
rect 25976 56 26004 1414
rect 26160 513 26188 2586
rect 26240 2576 26292 2582
rect 26240 2518 26292 2524
rect 26146 504 26202 513
rect 26146 439 26202 448
rect 26252 56 26280 2518
rect 26436 270 26464 3878
rect 26516 2304 26568 2310
rect 26516 2246 26568 2252
rect 26424 264 26476 270
rect 26424 206 26476 212
rect 26528 56 26556 2246
rect 26620 1290 26648 7278
rect 27010 6556 27318 6565
rect 27010 6554 27016 6556
rect 27072 6554 27096 6556
rect 27152 6554 27176 6556
rect 27232 6554 27256 6556
rect 27312 6554 27318 6556
rect 27072 6502 27074 6554
rect 27254 6502 27256 6554
rect 27010 6500 27016 6502
rect 27072 6500 27096 6502
rect 27152 6500 27176 6502
rect 27232 6500 27256 6502
rect 27312 6500 27318 6502
rect 27010 6491 27318 6500
rect 27010 5468 27318 5477
rect 27010 5466 27016 5468
rect 27072 5466 27096 5468
rect 27152 5466 27176 5468
rect 27232 5466 27256 5468
rect 27312 5466 27318 5468
rect 27072 5414 27074 5466
rect 27254 5414 27256 5466
rect 27010 5412 27016 5414
rect 27072 5412 27096 5414
rect 27152 5412 27176 5414
rect 27232 5412 27256 5414
rect 27312 5412 27318 5414
rect 27010 5403 27318 5412
rect 27632 4826 27660 8434
rect 28816 8424 28868 8430
rect 28816 8366 28868 8372
rect 27896 5160 27948 5166
rect 27896 5102 27948 5108
rect 27528 4820 27580 4826
rect 27528 4762 27580 4768
rect 27620 4820 27672 4826
rect 27620 4762 27672 4768
rect 27540 4570 27568 4762
rect 27540 4554 27844 4570
rect 27540 4548 27856 4554
rect 27540 4542 27804 4548
rect 27804 4490 27856 4496
rect 27908 4486 27936 5102
rect 28172 5024 28224 5030
rect 28172 4966 28224 4972
rect 28184 4486 28212 4966
rect 28828 4486 28856 8366
rect 30564 5024 30616 5030
rect 30564 4966 30616 4972
rect 29000 4616 29052 4622
rect 29000 4558 29052 4564
rect 27896 4480 27948 4486
rect 27896 4422 27948 4428
rect 28172 4480 28224 4486
rect 28172 4422 28224 4428
rect 28816 4480 28868 4486
rect 28816 4422 28868 4428
rect 27010 4380 27318 4389
rect 27010 4378 27016 4380
rect 27072 4378 27096 4380
rect 27152 4378 27176 4380
rect 27232 4378 27256 4380
rect 27312 4378 27318 4380
rect 27072 4326 27074 4378
rect 27254 4326 27256 4378
rect 27010 4324 27016 4326
rect 27072 4324 27096 4326
rect 27152 4324 27176 4326
rect 27232 4324 27256 4326
rect 27312 4324 27318 4326
rect 27010 4315 27318 4324
rect 29012 4214 29040 4558
rect 29000 4208 29052 4214
rect 29000 4150 29052 4156
rect 29644 4208 29696 4214
rect 29644 4150 29696 4156
rect 27804 4140 27856 4146
rect 27804 4082 27856 4088
rect 28356 4140 28408 4146
rect 28356 4082 28408 4088
rect 29184 4140 29236 4146
rect 29184 4082 29236 4088
rect 26700 3936 26752 3942
rect 26700 3878 26752 3884
rect 27436 3936 27488 3942
rect 27436 3878 27488 3884
rect 26712 2990 26740 3878
rect 27010 3292 27318 3301
rect 27010 3290 27016 3292
rect 27072 3290 27096 3292
rect 27152 3290 27176 3292
rect 27232 3290 27256 3292
rect 27312 3290 27318 3292
rect 27072 3238 27074 3290
rect 27254 3238 27256 3290
rect 27010 3236 27016 3238
rect 27072 3236 27096 3238
rect 27152 3236 27176 3238
rect 27232 3236 27256 3238
rect 27312 3236 27318 3238
rect 27010 3227 27318 3236
rect 27068 3188 27120 3194
rect 27068 3130 27120 3136
rect 26700 2984 26752 2990
rect 26700 2926 26752 2932
rect 26884 2848 26936 2854
rect 26884 2790 26936 2796
rect 26792 2644 26844 2650
rect 26792 2586 26844 2592
rect 26608 1284 26660 1290
rect 26608 1226 26660 1232
rect 26804 56 26832 2586
rect 15304 14 15424 42
rect 15474 0 15530 56
rect 15750 0 15806 56
rect 16026 0 16082 56
rect 16302 0 16358 56
rect 16578 0 16634 56
rect 16854 0 16910 56
rect 17130 0 17186 56
rect 17406 0 17462 56
rect 17682 0 17738 56
rect 17958 0 18014 56
rect 18234 0 18290 56
rect 18510 0 18566 56
rect 18786 0 18842 56
rect 19062 0 19118 56
rect 19338 0 19394 56
rect 19614 0 19670 56
rect 19890 0 19946 56
rect 20166 0 20222 56
rect 20442 0 20498 56
rect 20718 0 20774 56
rect 20994 0 21050 56
rect 21270 0 21326 56
rect 21546 0 21602 56
rect 21822 0 21878 56
rect 22098 0 22154 56
rect 22374 0 22430 56
rect 22650 0 22706 56
rect 22926 0 22982 56
rect 23202 0 23258 56
rect 23478 0 23534 56
rect 23754 0 23810 56
rect 24030 0 24086 56
rect 24306 0 24362 56
rect 24582 0 24638 56
rect 24858 0 24914 56
rect 25134 0 25190 56
rect 25410 0 25466 56
rect 25686 0 25742 56
rect 25962 0 26018 56
rect 26238 0 26294 56
rect 26514 0 26570 56
rect 26790 0 26846 56
rect 26896 42 26924 2790
rect 27080 2446 27108 3130
rect 27448 3058 27476 3878
rect 27436 3052 27488 3058
rect 27436 2994 27488 3000
rect 27344 2576 27396 2582
rect 27344 2518 27396 2524
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 27010 2204 27318 2213
rect 27010 2202 27016 2204
rect 27072 2202 27096 2204
rect 27152 2202 27176 2204
rect 27232 2202 27256 2204
rect 27312 2202 27318 2204
rect 27072 2150 27074 2202
rect 27254 2150 27256 2202
rect 27010 2148 27016 2150
rect 27072 2148 27096 2150
rect 27152 2148 27176 2150
rect 27232 2148 27256 2150
rect 27312 2148 27318 2150
rect 27010 2139 27318 2148
rect 26988 56 27108 82
rect 27356 56 27384 2518
rect 27712 2440 27764 2446
rect 27712 2382 27764 2388
rect 27620 2372 27672 2378
rect 27620 2314 27672 2320
rect 27632 56 27660 2314
rect 27724 1630 27752 2382
rect 27712 1624 27764 1630
rect 27712 1566 27764 1572
rect 27816 338 27844 4082
rect 28264 4004 28316 4010
rect 28264 3946 28316 3952
rect 27896 3936 27948 3942
rect 27896 3878 27948 3884
rect 27908 2446 27936 3878
rect 28172 2848 28224 2854
rect 28172 2790 28224 2796
rect 27988 2644 28040 2650
rect 27988 2586 28040 2592
rect 27896 2440 27948 2446
rect 27896 2382 27948 2388
rect 28000 1170 28028 2586
rect 27908 1142 28028 1170
rect 27804 332 27856 338
rect 27804 274 27856 280
rect 27908 56 27936 1142
rect 28184 56 28212 2790
rect 28276 1873 28304 3946
rect 28262 1864 28318 1873
rect 28262 1799 28318 1808
rect 28368 202 28396 4082
rect 28540 4072 28592 4078
rect 28540 4014 28592 4020
rect 28448 2848 28500 2854
rect 28448 2790 28500 2796
rect 28356 196 28408 202
rect 28356 138 28408 144
rect 28460 56 28488 2790
rect 28552 1766 28580 4014
rect 28632 3936 28684 3942
rect 28816 3936 28868 3942
rect 28684 3884 28764 3890
rect 28632 3878 28764 3884
rect 28816 3878 28868 3884
rect 28644 3862 28764 3878
rect 28736 3738 28764 3862
rect 28632 3732 28684 3738
rect 28632 3674 28684 3680
rect 28724 3732 28776 3738
rect 28724 3674 28776 3680
rect 28644 1834 28672 3674
rect 28724 2576 28776 2582
rect 28724 2518 28776 2524
rect 28632 1828 28684 1834
rect 28632 1770 28684 1776
rect 28540 1760 28592 1766
rect 28540 1702 28592 1708
rect 28736 56 28764 2518
rect 28828 2446 28856 3878
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 28920 2446 28948 3334
rect 28816 2440 28868 2446
rect 28816 2382 28868 2388
rect 28908 2440 28960 2446
rect 28908 2382 28960 2388
rect 29000 2304 29052 2310
rect 29000 2246 29052 2252
rect 29012 56 29040 2246
rect 29196 134 29224 4082
rect 29552 4072 29604 4078
rect 29380 4020 29552 4026
rect 29380 4014 29604 4020
rect 29380 3998 29592 4014
rect 29276 3528 29328 3534
rect 29274 3496 29276 3505
rect 29328 3496 29330 3505
rect 29274 3431 29330 3440
rect 29276 2848 29328 2854
rect 29276 2790 29328 2796
rect 29184 128 29236 134
rect 29184 70 29236 76
rect 29288 56 29316 2790
rect 29380 241 29408 3998
rect 29460 3936 29512 3942
rect 29460 3878 29512 3884
rect 29366 232 29422 241
rect 29366 167 29422 176
rect 29472 66 29500 3878
rect 29656 3618 29684 4150
rect 30288 4072 30340 4078
rect 29932 4020 30288 4026
rect 29932 4014 30340 4020
rect 29932 3998 30328 4014
rect 30472 4004 30524 4010
rect 29656 3590 29776 3618
rect 29644 3460 29696 3466
rect 29644 3402 29696 3408
rect 29552 3392 29604 3398
rect 29552 3334 29604 3340
rect 29564 3194 29592 3334
rect 29656 3194 29684 3402
rect 29552 3188 29604 3194
rect 29552 3130 29604 3136
rect 29644 3188 29696 3194
rect 29644 3130 29696 3136
rect 29748 3074 29776 3590
rect 29828 3392 29880 3398
rect 29828 3334 29880 3340
rect 29840 3126 29868 3334
rect 29656 3046 29776 3074
rect 29828 3120 29880 3126
rect 29828 3062 29880 3068
rect 29552 2100 29604 2106
rect 29552 2042 29604 2048
rect 29460 60 29512 66
rect 26988 54 27122 56
rect 26988 42 27016 54
rect 26896 14 27016 42
rect 27066 0 27122 54
rect 27342 0 27398 56
rect 27618 0 27674 56
rect 27894 0 27950 56
rect 28170 0 28226 56
rect 28446 0 28502 56
rect 28722 0 28778 56
rect 28998 0 29054 56
rect 29274 0 29330 56
rect 29564 56 29592 2042
rect 29656 1358 29684 3046
rect 29932 2774 29960 3998
rect 30472 3946 30524 3952
rect 30012 3936 30064 3942
rect 30012 3878 30064 3884
rect 30196 3936 30248 3942
rect 30196 3878 30248 3884
rect 30380 3936 30432 3942
rect 30380 3878 30432 3884
rect 29748 2746 29960 2774
rect 29748 2417 29776 2746
rect 29828 2644 29880 2650
rect 29828 2586 29880 2592
rect 29734 2408 29790 2417
rect 29734 2343 29790 2352
rect 29644 1352 29696 1358
rect 29644 1294 29696 1300
rect 29840 56 29868 2586
rect 30024 2514 30052 3878
rect 30104 2576 30156 2582
rect 30104 2518 30156 2524
rect 30012 2508 30064 2514
rect 30012 2450 30064 2456
rect 30116 56 30144 2518
rect 30208 2446 30236 3878
rect 30288 3392 30340 3398
rect 30288 3334 30340 3340
rect 30196 2440 30248 2446
rect 30196 2382 30248 2388
rect 30300 1902 30328 3334
rect 30392 3058 30420 3878
rect 30380 3052 30432 3058
rect 30380 2994 30432 3000
rect 30380 2848 30432 2854
rect 30380 2790 30432 2796
rect 30288 1896 30340 1902
rect 30288 1838 30340 1844
rect 30392 56 30420 2790
rect 30484 2774 30512 3946
rect 30576 3058 30604 4966
rect 30760 4826 30788 8434
rect 31312 5370 31340 8434
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 33010 7644 33318 7653
rect 33010 7642 33016 7644
rect 33072 7642 33096 7644
rect 33152 7642 33176 7644
rect 33232 7642 33256 7644
rect 33312 7642 33318 7644
rect 33072 7590 33074 7642
rect 33254 7590 33256 7642
rect 33010 7588 33016 7590
rect 33072 7588 33096 7590
rect 33152 7588 33176 7590
rect 33232 7588 33256 7590
rect 33312 7588 33318 7590
rect 33010 7579 33318 7588
rect 32588 7540 32640 7546
rect 32588 7482 32640 7488
rect 31852 7336 31904 7342
rect 31852 7278 31904 7284
rect 31758 6216 31814 6225
rect 31758 6151 31814 6160
rect 31116 5364 31168 5370
rect 31116 5306 31168 5312
rect 31300 5364 31352 5370
rect 31300 5306 31352 5312
rect 30748 4820 30800 4826
rect 30748 4762 30800 4768
rect 30840 4820 30892 4826
rect 30840 4762 30892 4768
rect 30852 4622 30880 4762
rect 31128 4758 31156 5306
rect 31392 5160 31444 5166
rect 31392 5102 31444 5108
rect 31116 4752 31168 4758
rect 31116 4694 31168 4700
rect 30840 4616 30892 4622
rect 30840 4558 30892 4564
rect 31300 4072 31352 4078
rect 31300 4014 31352 4020
rect 30840 3936 30892 3942
rect 30840 3878 30892 3884
rect 31116 3936 31168 3942
rect 31116 3878 31168 3884
rect 30564 3052 30616 3058
rect 30564 2994 30616 3000
rect 30484 2746 30604 2774
rect 30472 2576 30524 2582
rect 30472 2518 30524 2524
rect 30484 2106 30512 2518
rect 30576 2446 30604 2746
rect 30656 2576 30708 2582
rect 30656 2518 30708 2524
rect 30564 2440 30616 2446
rect 30564 2382 30616 2388
rect 30472 2100 30524 2106
rect 30472 2042 30524 2048
rect 30472 1896 30524 1902
rect 30472 1838 30524 1844
rect 30484 1562 30512 1838
rect 30472 1556 30524 1562
rect 30472 1498 30524 1504
rect 30668 56 30696 2518
rect 30852 105 30880 3878
rect 31024 3732 31076 3738
rect 31024 3674 31076 3680
rect 30932 2848 30984 2854
rect 30932 2790 30984 2796
rect 30838 96 30894 105
rect 29460 2 29512 8
rect 29550 0 29606 56
rect 29826 0 29882 56
rect 30102 0 30158 56
rect 30378 0 30434 56
rect 30654 0 30710 56
rect 30944 56 30972 2790
rect 31036 2446 31064 3674
rect 31024 2440 31076 2446
rect 31024 2382 31076 2388
rect 31128 2310 31156 3878
rect 31312 2922 31340 4014
rect 31300 2916 31352 2922
rect 31300 2858 31352 2864
rect 31404 2446 31432 5102
rect 31392 2440 31444 2446
rect 31392 2382 31444 2388
rect 31116 2304 31168 2310
rect 31116 2246 31168 2252
rect 31300 2304 31352 2310
rect 31300 2246 31352 2252
rect 31312 1170 31340 2246
rect 31482 1456 31538 1465
rect 31482 1391 31538 1400
rect 31220 1142 31340 1170
rect 31220 56 31248 1142
rect 31496 56 31524 1391
rect 31772 56 31800 6151
rect 30838 31 30894 40
rect 30930 0 30986 56
rect 31206 0 31262 56
rect 31482 0 31538 56
rect 31758 0 31814 56
rect 31864 42 31892 7278
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 32128 2440 32180 2446
rect 32128 2382 32180 2388
rect 32220 2440 32272 2446
rect 32220 2382 32272 2388
rect 32140 1834 32168 2382
rect 32232 2106 32260 2382
rect 32220 2100 32272 2106
rect 32220 2042 32272 2048
rect 32128 1828 32180 1834
rect 32128 1770 32180 1776
rect 32312 400 32364 406
rect 32312 342 32364 348
rect 31956 56 32076 82
rect 32324 56 32352 342
rect 32600 56 32628 7482
rect 33414 7440 33470 7449
rect 33414 7375 33470 7384
rect 33968 7404 34020 7410
rect 33010 6556 33318 6565
rect 33010 6554 33016 6556
rect 33072 6554 33096 6556
rect 33152 6554 33176 6556
rect 33232 6554 33256 6556
rect 33312 6554 33318 6556
rect 33072 6502 33074 6554
rect 33254 6502 33256 6554
rect 33010 6500 33016 6502
rect 33072 6500 33096 6502
rect 33152 6500 33176 6502
rect 33232 6500 33256 6502
rect 33312 6500 33318 6502
rect 33010 6491 33318 6500
rect 33010 5468 33318 5477
rect 33010 5466 33016 5468
rect 33072 5466 33096 5468
rect 33152 5466 33176 5468
rect 33232 5466 33256 5468
rect 33312 5466 33318 5468
rect 33072 5414 33074 5466
rect 33254 5414 33256 5466
rect 33010 5412 33016 5414
rect 33072 5412 33096 5414
rect 33152 5412 33176 5414
rect 33232 5412 33256 5414
rect 33312 5412 33318 5414
rect 33010 5403 33318 5412
rect 33010 4380 33318 4389
rect 33010 4378 33016 4380
rect 33072 4378 33096 4380
rect 33152 4378 33176 4380
rect 33232 4378 33256 4380
rect 33312 4378 33318 4380
rect 33072 4326 33074 4378
rect 33254 4326 33256 4378
rect 33010 4324 33016 4326
rect 33072 4324 33096 4326
rect 33152 4324 33176 4326
rect 33232 4324 33256 4326
rect 33312 4324 33318 4326
rect 33010 4315 33318 4324
rect 33010 3292 33318 3301
rect 33010 3290 33016 3292
rect 33072 3290 33096 3292
rect 33152 3290 33176 3292
rect 33232 3290 33256 3292
rect 33312 3290 33318 3292
rect 33072 3238 33074 3290
rect 33254 3238 33256 3290
rect 33010 3236 33016 3238
rect 33072 3236 33096 3238
rect 33152 3236 33176 3238
rect 33232 3236 33256 3238
rect 33312 3236 33318 3238
rect 33010 3227 33318 3236
rect 33138 2952 33194 2961
rect 33138 2887 33194 2896
rect 32862 2544 32918 2553
rect 33152 2514 33180 2887
rect 32862 2479 32918 2488
rect 33140 2508 33192 2514
rect 32876 56 32904 2479
rect 33140 2450 33192 2456
rect 33010 2204 33318 2213
rect 33010 2202 33016 2204
rect 33072 2202 33096 2204
rect 33152 2202 33176 2204
rect 33232 2202 33256 2204
rect 33312 2202 33318 2204
rect 33072 2150 33074 2202
rect 33254 2150 33256 2202
rect 33010 2148 33016 2150
rect 33072 2148 33096 2150
rect 33152 2148 33176 2150
rect 33232 2148 33256 2150
rect 33312 2148 33318 2150
rect 33010 2139 33318 2148
rect 33428 218 33456 7375
rect 33968 7346 34020 7352
rect 33506 3632 33562 3641
rect 33506 3567 33562 3576
rect 33520 2582 33548 3567
rect 33508 2576 33560 2582
rect 33508 2518 33560 2524
rect 33692 1284 33744 1290
rect 33692 1226 33744 1232
rect 33508 468 33560 474
rect 33508 410 33560 416
rect 33336 190 33456 218
rect 33152 56 33272 82
rect 31956 54 32090 56
rect 31956 42 31984 54
rect 31864 14 31984 42
rect 32034 0 32090 54
rect 32310 0 32366 56
rect 32586 0 32642 56
rect 32862 0 32918 56
rect 33138 54 33272 56
rect 33138 0 33194 54
rect 33244 42 33272 54
rect 33336 42 33364 190
rect 33520 82 33548 410
rect 33428 56 33548 82
rect 33704 56 33732 1226
rect 33980 56 34008 7346
rect 34152 6792 34204 6798
rect 34152 6734 34204 6740
rect 34164 2774 34192 6734
rect 34256 5914 34284 8434
rect 34992 5914 35020 8434
rect 36832 5914 36860 8434
rect 36924 8090 36952 9279
rect 37278 9072 37334 9081
rect 37278 9007 37334 9016
rect 37292 8090 37320 9007
rect 37832 8968 37884 8974
rect 37832 8910 37884 8916
rect 37646 8528 37702 8537
rect 37844 8498 37872 8910
rect 38304 8634 38332 11096
rect 38474 8800 38530 8809
rect 38474 8735 38530 8744
rect 38292 8628 38344 8634
rect 38292 8570 38344 8576
rect 37646 8463 37702 8472
rect 37832 8492 37884 8498
rect 37556 8424 37608 8430
rect 37556 8366 37608 8372
rect 36912 8084 36964 8090
rect 36912 8026 36964 8032
rect 37280 8084 37332 8090
rect 37280 8026 37332 8032
rect 37096 7880 37148 7886
rect 37096 7822 37148 7828
rect 37464 7880 37516 7886
rect 37464 7822 37516 7828
rect 37108 7002 37136 7822
rect 37280 7336 37332 7342
rect 37280 7278 37332 7284
rect 37096 6996 37148 7002
rect 37096 6938 37148 6944
rect 37292 6458 37320 7278
rect 37476 7274 37504 7822
rect 37464 7268 37516 7274
rect 37464 7210 37516 7216
rect 37280 6452 37332 6458
rect 37280 6394 37332 6400
rect 37568 5914 37596 8366
rect 37660 8090 37688 8463
rect 37832 8434 37884 8440
rect 37950 8188 38258 8197
rect 37950 8186 37956 8188
rect 38012 8186 38036 8188
rect 38092 8186 38116 8188
rect 38172 8186 38196 8188
rect 38252 8186 38258 8188
rect 38012 8134 38014 8186
rect 38194 8134 38196 8186
rect 37950 8132 37956 8134
rect 38012 8132 38036 8134
rect 38092 8132 38116 8134
rect 38172 8132 38196 8134
rect 38252 8132 38258 8134
rect 37950 8123 38258 8132
rect 37648 8084 37700 8090
rect 37648 8026 37700 8032
rect 38016 7744 38068 7750
rect 38384 7744 38436 7750
rect 38016 7686 38068 7692
rect 38382 7712 38384 7721
rect 38436 7712 38438 7721
rect 38028 7449 38056 7686
rect 38382 7647 38438 7656
rect 38488 7546 38516 8735
rect 38936 8560 38988 8566
rect 38936 8502 38988 8508
rect 38752 8356 38804 8362
rect 38752 8298 38804 8304
rect 38764 8265 38792 8298
rect 38750 8256 38806 8265
rect 38750 8191 38806 8200
rect 38948 7993 38976 8502
rect 38934 7984 38990 7993
rect 38934 7919 38990 7928
rect 38476 7540 38528 7546
rect 38476 7482 38528 7488
rect 38014 7440 38070 7449
rect 38014 7375 38070 7384
rect 38384 7200 38436 7206
rect 38382 7168 38384 7177
rect 38436 7168 38438 7177
rect 37950 7100 38258 7109
rect 38382 7103 38438 7112
rect 37950 7098 37956 7100
rect 38012 7098 38036 7100
rect 38092 7098 38116 7100
rect 38172 7098 38196 7100
rect 38252 7098 38258 7100
rect 38012 7046 38014 7098
rect 38194 7046 38196 7098
rect 37950 7044 37956 7046
rect 38012 7044 38036 7046
rect 38092 7044 38116 7046
rect 38172 7044 38196 7046
rect 38252 7044 38258 7046
rect 37950 7035 38258 7044
rect 38198 6896 38254 6905
rect 38198 6831 38254 6840
rect 38382 6896 38438 6905
rect 38382 6831 38438 6840
rect 38212 6798 38240 6831
rect 38200 6792 38252 6798
rect 38200 6734 38252 6740
rect 38396 6662 38424 6831
rect 38016 6656 38068 6662
rect 38014 6624 38016 6633
rect 38384 6656 38436 6662
rect 38068 6624 38070 6633
rect 38384 6598 38436 6604
rect 38014 6559 38070 6568
rect 38384 6452 38436 6458
rect 38384 6394 38436 6400
rect 38396 6361 38424 6394
rect 38382 6352 38438 6361
rect 38382 6287 38438 6296
rect 37832 6180 37884 6186
rect 37832 6122 37884 6128
rect 34244 5908 34296 5914
rect 34244 5850 34296 5856
rect 34980 5908 35032 5914
rect 34980 5850 35032 5856
rect 36820 5908 36872 5914
rect 36820 5850 36872 5856
rect 37556 5908 37608 5914
rect 37556 5850 37608 5856
rect 34520 5840 34572 5846
rect 34520 5782 34572 5788
rect 34164 2746 34284 2774
rect 34256 56 34284 2746
rect 34532 56 34560 5782
rect 36176 5772 36228 5778
rect 36176 5714 36228 5720
rect 35992 5228 36044 5234
rect 35992 5170 36044 5176
rect 35348 4820 35400 4826
rect 35348 4762 35400 4768
rect 35072 1760 35124 1766
rect 35072 1702 35124 1708
rect 34796 1352 34848 1358
rect 34796 1294 34848 1300
rect 34808 56 34836 1294
rect 35084 56 35112 1702
rect 35360 56 35388 4762
rect 35624 4684 35676 4690
rect 35624 4626 35676 4632
rect 35636 56 35664 4626
rect 35898 4040 35954 4049
rect 35898 3975 35954 3984
rect 35912 3602 35940 3975
rect 35900 3596 35952 3602
rect 35900 3538 35952 3544
rect 36004 2774 36032 5170
rect 35912 2746 36032 2774
rect 35912 56 35940 2746
rect 36188 56 36216 5714
rect 37844 5710 37872 6122
rect 39120 6112 39172 6118
rect 39118 6080 39120 6089
rect 39172 6080 39174 6089
rect 37950 6012 38258 6021
rect 39118 6015 39174 6024
rect 37950 6010 37956 6012
rect 38012 6010 38036 6012
rect 38092 6010 38116 6012
rect 38172 6010 38196 6012
rect 38252 6010 38258 6012
rect 38012 5958 38014 6010
rect 38194 5958 38196 6010
rect 37950 5956 37956 5958
rect 38012 5956 38036 5958
rect 38092 5956 38116 5958
rect 38172 5956 38196 5958
rect 38252 5956 38258 5958
rect 37950 5947 38258 5956
rect 38384 5840 38436 5846
rect 38382 5808 38384 5817
rect 38436 5808 38438 5817
rect 38382 5743 38438 5752
rect 36452 5704 36504 5710
rect 36452 5646 36504 5652
rect 36728 5704 36780 5710
rect 36728 5646 36780 5652
rect 37004 5704 37056 5710
rect 37004 5646 37056 5652
rect 37832 5704 37884 5710
rect 37832 5646 37884 5652
rect 36464 56 36492 5646
rect 36636 2304 36688 2310
rect 36636 2246 36688 2252
rect 36648 2009 36676 2246
rect 36634 2000 36690 2009
rect 36634 1935 36690 1944
rect 36740 56 36768 5646
rect 36820 2440 36872 2446
rect 36820 2382 36872 2388
rect 36832 1902 36860 2382
rect 36820 1896 36872 1902
rect 36820 1838 36872 1844
rect 37016 56 37044 5646
rect 38016 5568 38068 5574
rect 38014 5536 38016 5545
rect 38068 5536 38070 5545
rect 38014 5471 38070 5480
rect 38384 5364 38436 5370
rect 38384 5306 38436 5312
rect 38396 5273 38424 5306
rect 38382 5264 38438 5273
rect 38382 5199 38438 5208
rect 39120 5024 39172 5030
rect 39118 4992 39120 5001
rect 39172 4992 39174 5001
rect 37950 4924 38258 4933
rect 39118 4927 39174 4936
rect 37950 4922 37956 4924
rect 38012 4922 38036 4924
rect 38092 4922 38116 4924
rect 38172 4922 38196 4924
rect 38252 4922 38258 4924
rect 38012 4870 38014 4922
rect 38194 4870 38196 4922
rect 37950 4868 37956 4870
rect 38012 4868 38036 4870
rect 38092 4868 38116 4870
rect 38172 4868 38196 4870
rect 38252 4868 38258 4870
rect 37950 4859 38258 4868
rect 38200 4752 38252 4758
rect 38384 4752 38436 4758
rect 38200 4694 38252 4700
rect 38382 4720 38384 4729
rect 38436 4720 38438 4729
rect 38016 4480 38068 4486
rect 38014 4448 38016 4457
rect 38068 4448 38070 4457
rect 38014 4383 38070 4392
rect 38212 4146 38240 4694
rect 38382 4655 38438 4664
rect 38382 4176 38438 4185
rect 38200 4140 38252 4146
rect 38382 4111 38438 4120
rect 38200 4082 38252 4088
rect 37464 4072 37516 4078
rect 37464 4014 37516 4020
rect 37476 3058 37504 4014
rect 38396 4010 38424 4111
rect 38384 4004 38436 4010
rect 38384 3946 38436 3952
rect 39120 3936 39172 3942
rect 39118 3904 39120 3913
rect 39172 3904 39174 3913
rect 37950 3836 38258 3845
rect 39118 3839 39174 3848
rect 37950 3834 37956 3836
rect 38012 3834 38036 3836
rect 38092 3834 38116 3836
rect 38172 3834 38196 3836
rect 38252 3834 38258 3836
rect 38012 3782 38014 3834
rect 38194 3782 38196 3834
rect 37950 3780 37956 3782
rect 38012 3780 38036 3782
rect 38092 3780 38116 3782
rect 38172 3780 38196 3782
rect 38252 3780 38258 3782
rect 37950 3771 38258 3780
rect 38384 3664 38436 3670
rect 38382 3632 38384 3641
rect 38436 3632 38438 3641
rect 38382 3567 38438 3576
rect 37924 3460 37976 3466
rect 37924 3402 37976 3408
rect 37936 3058 37964 3402
rect 38016 3392 38068 3398
rect 38014 3360 38016 3369
rect 38068 3360 38070 3369
rect 38014 3295 38070 3304
rect 38384 3188 38436 3194
rect 38384 3130 38436 3136
rect 38396 3097 38424 3130
rect 38382 3088 38438 3097
rect 37464 3052 37516 3058
rect 37464 2994 37516 3000
rect 37924 3052 37976 3058
rect 38382 3023 38438 3032
rect 37924 2994 37976 3000
rect 37832 2848 37884 2854
rect 39120 2848 39172 2854
rect 37832 2790 37884 2796
rect 39118 2816 39120 2825
rect 39172 2816 39174 2825
rect 37188 2304 37240 2310
rect 37188 2246 37240 2252
rect 37648 2304 37700 2310
rect 37648 2246 37700 2252
rect 37200 1465 37228 2246
rect 37186 1456 37242 1465
rect 37186 1391 37242 1400
rect 37660 1193 37688 2246
rect 37844 1737 37872 2790
rect 37950 2748 38258 2757
rect 39118 2751 39174 2760
rect 37950 2746 37956 2748
rect 38012 2746 38036 2748
rect 38092 2746 38116 2748
rect 38172 2746 38196 2748
rect 38252 2746 38258 2748
rect 38012 2694 38014 2746
rect 38194 2694 38196 2746
rect 37950 2692 37956 2694
rect 38012 2692 38036 2694
rect 38092 2692 38116 2694
rect 38172 2692 38196 2694
rect 38252 2692 38258 2694
rect 37950 2683 38258 2692
rect 38384 2576 38436 2582
rect 38382 2544 38384 2553
rect 38436 2544 38438 2553
rect 38382 2479 38438 2488
rect 38200 2440 38252 2446
rect 38200 2382 38252 2388
rect 38016 2304 38068 2310
rect 38014 2272 38016 2281
rect 38068 2272 38070 2281
rect 38014 2207 38070 2216
rect 38212 2038 38240 2382
rect 38200 2032 38252 2038
rect 38200 1974 38252 1980
rect 37830 1728 37886 1737
rect 37830 1663 37886 1672
rect 37646 1184 37702 1193
rect 37646 1119 37702 1128
rect 33244 14 33364 42
rect 33414 54 33548 56
rect 33414 0 33470 54
rect 33690 0 33746 56
rect 33966 0 34022 56
rect 34242 0 34298 56
rect 34518 0 34574 56
rect 34794 0 34850 56
rect 35070 0 35126 56
rect 35346 0 35402 56
rect 35622 0 35678 56
rect 35898 0 35954 56
rect 36174 0 36230 56
rect 36450 0 36506 56
rect 36726 0 36782 56
rect 37002 0 37058 56
<< via2 >>
rect 2870 8744 2926 8800
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 9176 8730 9232 8732
rect 9256 8730 9312 8732
rect 9016 8678 9062 8730
rect 9062 8678 9072 8730
rect 9096 8678 9126 8730
rect 9126 8678 9138 8730
rect 9138 8678 9152 8730
rect 9176 8678 9190 8730
rect 9190 8678 9202 8730
rect 9202 8678 9232 8730
rect 9256 8678 9266 8730
rect 9266 8678 9312 8730
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 9176 8676 9232 8678
rect 9256 8676 9312 8678
rect 14646 9288 14702 9344
rect 2870 8336 2926 8392
rect 1766 8200 1822 8256
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 13956 8186 14012 8188
rect 14036 8186 14092 8188
rect 14116 8186 14172 8188
rect 14196 8186 14252 8188
rect 13956 8134 14002 8186
rect 14002 8134 14012 8186
rect 14036 8134 14066 8186
rect 14066 8134 14078 8186
rect 14078 8134 14092 8186
rect 14116 8134 14130 8186
rect 14130 8134 14142 8186
rect 14142 8134 14172 8186
rect 14196 8134 14206 8186
rect 14206 8134 14252 8186
rect 13956 8132 14012 8134
rect 14036 8132 14092 8134
rect 14116 8132 14172 8134
rect 14196 8132 14252 8134
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 9176 7642 9232 7644
rect 9256 7642 9312 7644
rect 9016 7590 9062 7642
rect 9062 7590 9072 7642
rect 9096 7590 9126 7642
rect 9126 7590 9138 7642
rect 9138 7590 9152 7642
rect 9176 7590 9190 7642
rect 9190 7590 9202 7642
rect 9202 7590 9232 7642
rect 9256 7590 9266 7642
rect 9266 7590 9312 7642
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 9176 7588 9232 7590
rect 9256 7588 9312 7590
rect 14830 9016 14886 9072
rect 15016 8730 15072 8732
rect 15096 8730 15152 8732
rect 15176 8730 15232 8732
rect 15256 8730 15312 8732
rect 15016 8678 15062 8730
rect 15062 8678 15072 8730
rect 15096 8678 15126 8730
rect 15126 8678 15138 8730
rect 15138 8678 15152 8730
rect 15176 8678 15190 8730
rect 15190 8678 15202 8730
rect 15202 8678 15232 8730
rect 15256 8678 15266 8730
rect 15266 8678 15312 8730
rect 15016 8676 15072 8678
rect 15096 8676 15152 8678
rect 15176 8676 15232 8678
rect 15256 8676 15312 8678
rect 14922 8336 14978 8392
rect 15016 7642 15072 7644
rect 15096 7642 15152 7644
rect 15176 7642 15232 7644
rect 15256 7642 15312 7644
rect 15016 7590 15062 7642
rect 15062 7590 15072 7642
rect 15096 7590 15126 7642
rect 15126 7590 15138 7642
rect 15138 7590 15152 7642
rect 15176 7590 15190 7642
rect 15190 7590 15202 7642
rect 15202 7590 15232 7642
rect 15256 7590 15266 7642
rect 15266 7590 15312 7642
rect 15016 7588 15072 7590
rect 15096 7588 15152 7590
rect 15176 7588 15232 7590
rect 15256 7588 15312 7590
rect 15290 7404 15346 7440
rect 15290 7384 15292 7404
rect 15292 7384 15344 7404
rect 15344 7384 15346 7404
rect 1766 7248 1822 7304
rect 19798 9560 19854 9616
rect 17038 8472 17094 8528
rect 18234 7928 18290 7984
rect 18050 7792 18106 7848
rect 18602 7792 18658 7848
rect 19522 7248 19578 7304
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 20196 8186 20252 8188
rect 19956 8134 20002 8186
rect 20002 8134 20012 8186
rect 20036 8134 20066 8186
rect 20066 8134 20078 8186
rect 20078 8134 20092 8186
rect 20116 8134 20130 8186
rect 20130 8134 20142 8186
rect 20142 8134 20172 8186
rect 20196 8134 20206 8186
rect 20206 8134 20252 8186
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 20196 8132 20252 8134
rect 20258 7248 20314 7304
rect 21016 8730 21072 8732
rect 21096 8730 21152 8732
rect 21176 8730 21232 8732
rect 21256 8730 21312 8732
rect 21016 8678 21062 8730
rect 21062 8678 21072 8730
rect 21096 8678 21126 8730
rect 21126 8678 21138 8730
rect 21138 8678 21152 8730
rect 21176 8678 21190 8730
rect 21190 8678 21202 8730
rect 21202 8678 21232 8730
rect 21256 8678 21266 8730
rect 21266 8678 21312 8730
rect 21016 8676 21072 8678
rect 21096 8676 21152 8678
rect 21176 8676 21232 8678
rect 21256 8676 21312 8678
rect 21016 7642 21072 7644
rect 21096 7642 21152 7644
rect 21176 7642 21232 7644
rect 21256 7642 21312 7644
rect 21016 7590 21062 7642
rect 21062 7590 21072 7642
rect 21096 7590 21126 7642
rect 21126 7590 21138 7642
rect 21138 7590 21152 7642
rect 21176 7590 21190 7642
rect 21190 7590 21202 7642
rect 21202 7590 21232 7642
rect 21256 7590 21266 7642
rect 21266 7590 21312 7642
rect 21016 7588 21072 7590
rect 21096 7588 21152 7590
rect 21176 7588 21232 7590
rect 21256 7588 21312 7590
rect 1306 7112 1362 7168
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 13956 7098 14012 7100
rect 14036 7098 14092 7100
rect 14116 7098 14172 7100
rect 14196 7098 14252 7100
rect 13956 7046 14002 7098
rect 14002 7046 14012 7098
rect 14036 7046 14066 7098
rect 14066 7046 14078 7098
rect 14078 7046 14092 7098
rect 14116 7046 14130 7098
rect 14130 7046 14142 7098
rect 14142 7046 14172 7098
rect 14196 7046 14206 7098
rect 14206 7046 14252 7098
rect 13956 7044 14012 7046
rect 14036 7044 14092 7046
rect 14116 7044 14172 7046
rect 14196 7044 14252 7046
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 20196 7098 20252 7100
rect 19956 7046 20002 7098
rect 20002 7046 20012 7098
rect 20036 7046 20066 7098
rect 20066 7046 20078 7098
rect 20078 7046 20092 7098
rect 20116 7046 20130 7098
rect 20130 7046 20142 7098
rect 20142 7046 20172 7098
rect 20196 7046 20206 7098
rect 20206 7046 20252 7098
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 20196 7044 20252 7046
rect 15750 6860 15806 6896
rect 15750 6840 15752 6860
rect 15752 6840 15804 6860
rect 15804 6840 15806 6860
rect 16118 6840 16174 6896
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 3882 5616 3938 5672
rect 2870 5480 2926 5536
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 2778 5208 2834 5264
rect 2962 5208 3018 5264
rect 2962 5072 3018 5128
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 570 2488 626 2544
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 4434 4392 4490 4448
rect 5722 1944 5778 2000
rect 5630 1400 5686 1456
rect 7654 4936 7710 4992
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 8298 5616 8354 5672
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 8390 4392 8446 4448
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 9176 6554 9232 6556
rect 9256 6554 9312 6556
rect 9016 6502 9062 6554
rect 9062 6502 9072 6554
rect 9096 6502 9126 6554
rect 9126 6502 9138 6554
rect 9138 6502 9152 6554
rect 9176 6502 9190 6554
rect 9190 6502 9202 6554
rect 9202 6502 9232 6554
rect 9256 6502 9266 6554
rect 9266 6502 9312 6554
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 9176 6500 9232 6502
rect 9256 6500 9312 6502
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 9176 5466 9232 5468
rect 9256 5466 9312 5468
rect 9016 5414 9062 5466
rect 9062 5414 9072 5466
rect 9096 5414 9126 5466
rect 9126 5414 9138 5466
rect 9138 5414 9152 5466
rect 9176 5414 9190 5466
rect 9190 5414 9202 5466
rect 9202 5414 9232 5466
rect 9256 5414 9266 5466
rect 9266 5414 9312 5466
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 9176 5412 9232 5414
rect 9256 5412 9312 5414
rect 9954 5616 10010 5672
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 9176 4378 9232 4380
rect 9256 4378 9312 4380
rect 9016 4326 9062 4378
rect 9062 4326 9072 4378
rect 9096 4326 9126 4378
rect 9126 4326 9138 4378
rect 9138 4326 9152 4378
rect 9176 4326 9190 4378
rect 9190 4326 9202 4378
rect 9202 4326 9232 4378
rect 9256 4326 9266 4378
rect 9266 4326 9312 4378
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 9176 4324 9232 4326
rect 9256 4324 9312 4326
rect 8758 3848 8814 3904
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 9176 3290 9232 3292
rect 9256 3290 9312 3292
rect 9016 3238 9062 3290
rect 9062 3238 9072 3290
rect 9096 3238 9126 3290
rect 9126 3238 9138 3290
rect 9138 3238 9152 3290
rect 9176 3238 9190 3290
rect 9190 3238 9202 3290
rect 9202 3238 9232 3290
rect 9256 3238 9266 3290
rect 9266 3238 9312 3290
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 9176 3236 9232 3238
rect 9256 3236 9312 3238
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 9176 2202 9232 2204
rect 9256 2202 9312 2204
rect 9016 2150 9062 2202
rect 9062 2150 9072 2202
rect 9096 2150 9126 2202
rect 9126 2150 9138 2202
rect 9138 2150 9152 2202
rect 9176 2150 9190 2202
rect 9190 2150 9202 2202
rect 9202 2150 9232 2202
rect 9256 2150 9266 2202
rect 9266 2150 9312 2202
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 9176 2148 9232 2150
rect 9256 2148 9312 2150
rect 9586 1672 9642 1728
rect 9954 1944 10010 2000
rect 11058 3984 11114 4040
rect 10966 2352 11022 2408
rect 11150 3168 11206 3224
rect 11242 2352 11298 2408
rect 11150 1536 11206 1592
rect 11610 2624 11666 2680
rect 16670 6704 16726 6760
rect 15016 6554 15072 6556
rect 15096 6554 15152 6556
rect 15176 6554 15232 6556
rect 15256 6554 15312 6556
rect 15016 6502 15062 6554
rect 15062 6502 15072 6554
rect 15096 6502 15126 6554
rect 15126 6502 15138 6554
rect 15138 6502 15152 6554
rect 15176 6502 15190 6554
rect 15190 6502 15202 6554
rect 15202 6502 15232 6554
rect 15256 6502 15266 6554
rect 15266 6502 15312 6554
rect 15016 6500 15072 6502
rect 15096 6500 15152 6502
rect 15176 6500 15232 6502
rect 15256 6500 15312 6502
rect 21016 6554 21072 6556
rect 21096 6554 21152 6556
rect 21176 6554 21232 6556
rect 21256 6554 21312 6556
rect 21016 6502 21062 6554
rect 21062 6502 21072 6554
rect 21096 6502 21126 6554
rect 21126 6502 21138 6554
rect 21138 6502 21152 6554
rect 21176 6502 21190 6554
rect 21190 6502 21202 6554
rect 21202 6502 21232 6554
rect 21256 6502 21266 6554
rect 21266 6502 21312 6554
rect 21016 6500 21072 6502
rect 21096 6500 21152 6502
rect 21176 6500 21232 6502
rect 21256 6500 21312 6502
rect 11886 2488 11942 2544
rect 13956 6010 14012 6012
rect 14036 6010 14092 6012
rect 14116 6010 14172 6012
rect 14196 6010 14252 6012
rect 13956 5958 14002 6010
rect 14002 5958 14012 6010
rect 14036 5958 14066 6010
rect 14066 5958 14078 6010
rect 14078 5958 14092 6010
rect 14116 5958 14130 6010
rect 14130 5958 14142 6010
rect 14142 5958 14172 6010
rect 14196 5958 14206 6010
rect 14206 5958 14252 6010
rect 13956 5956 14012 5958
rect 14036 5956 14092 5958
rect 14116 5956 14172 5958
rect 14196 5956 14252 5958
rect 18694 6296 18750 6352
rect 13174 2624 13230 2680
rect 13956 4922 14012 4924
rect 14036 4922 14092 4924
rect 14116 4922 14172 4924
rect 14196 4922 14252 4924
rect 13956 4870 14002 4922
rect 14002 4870 14012 4922
rect 14036 4870 14066 4922
rect 14066 4870 14078 4922
rect 14078 4870 14092 4922
rect 14116 4870 14130 4922
rect 14130 4870 14142 4922
rect 14142 4870 14172 4922
rect 14196 4870 14206 4922
rect 14206 4870 14252 4922
rect 13956 4868 14012 4870
rect 14036 4868 14092 4870
rect 14116 4868 14172 4870
rect 14196 4868 14252 4870
rect 13542 2488 13598 2544
rect 13956 3834 14012 3836
rect 14036 3834 14092 3836
rect 14116 3834 14172 3836
rect 14196 3834 14252 3836
rect 13956 3782 14002 3834
rect 14002 3782 14012 3834
rect 14036 3782 14066 3834
rect 14066 3782 14078 3834
rect 14078 3782 14092 3834
rect 14116 3782 14130 3834
rect 14130 3782 14142 3834
rect 14142 3782 14172 3834
rect 14196 3782 14206 3834
rect 14206 3782 14252 3834
rect 13956 3780 14012 3782
rect 14036 3780 14092 3782
rect 14116 3780 14172 3782
rect 14196 3780 14252 3782
rect 13956 2746 14012 2748
rect 14036 2746 14092 2748
rect 14116 2746 14172 2748
rect 14196 2746 14252 2748
rect 13956 2694 14002 2746
rect 14002 2694 14012 2746
rect 14036 2694 14066 2746
rect 14066 2694 14078 2746
rect 14078 2694 14092 2746
rect 14116 2694 14130 2746
rect 14130 2694 14142 2746
rect 14142 2694 14172 2746
rect 14196 2694 14206 2746
rect 14206 2694 14252 2746
rect 13956 2692 14012 2694
rect 14036 2692 14092 2694
rect 14116 2692 14172 2694
rect 14196 2692 14252 2694
rect 17406 6160 17462 6216
rect 15016 5466 15072 5468
rect 15096 5466 15152 5468
rect 15176 5466 15232 5468
rect 15256 5466 15312 5468
rect 15016 5414 15062 5466
rect 15062 5414 15072 5466
rect 15096 5414 15126 5466
rect 15126 5414 15138 5466
rect 15138 5414 15152 5466
rect 15176 5414 15190 5466
rect 15190 5414 15202 5466
rect 15202 5414 15232 5466
rect 15256 5414 15266 5466
rect 15266 5414 15312 5466
rect 15016 5412 15072 5414
rect 15096 5412 15152 5414
rect 15176 5412 15232 5414
rect 15256 5412 15312 5414
rect 15016 4378 15072 4380
rect 15096 4378 15152 4380
rect 15176 4378 15232 4380
rect 15256 4378 15312 4380
rect 15016 4326 15062 4378
rect 15062 4326 15072 4378
rect 15096 4326 15126 4378
rect 15126 4326 15138 4378
rect 15138 4326 15152 4378
rect 15176 4326 15190 4378
rect 15190 4326 15202 4378
rect 15202 4326 15232 4378
rect 15256 4326 15266 4378
rect 15266 4326 15312 4378
rect 15016 4324 15072 4326
rect 15096 4324 15152 4326
rect 15176 4324 15232 4326
rect 15256 4324 15312 4326
rect 15016 3290 15072 3292
rect 15096 3290 15152 3292
rect 15176 3290 15232 3292
rect 15256 3290 15312 3292
rect 15016 3238 15062 3290
rect 15062 3238 15072 3290
rect 15096 3238 15126 3290
rect 15126 3238 15138 3290
rect 15138 3238 15152 3290
rect 15176 3238 15190 3290
rect 15190 3238 15202 3290
rect 15202 3238 15232 3290
rect 15256 3238 15266 3290
rect 15266 3238 15312 3290
rect 15016 3236 15072 3238
rect 15096 3236 15152 3238
rect 15176 3236 15232 3238
rect 15256 3236 15312 3238
rect 15474 2352 15530 2408
rect 15016 2202 15072 2204
rect 15096 2202 15152 2204
rect 15176 2202 15232 2204
rect 15256 2202 15312 2204
rect 15016 2150 15062 2202
rect 15062 2150 15072 2202
rect 15096 2150 15126 2202
rect 15126 2150 15138 2202
rect 15138 2150 15152 2202
rect 15176 2150 15190 2202
rect 15190 2150 15202 2202
rect 15202 2150 15232 2202
rect 15256 2150 15266 2202
rect 15266 2150 15312 2202
rect 15016 2148 15072 2150
rect 15096 2148 15152 2150
rect 15176 2148 15232 2150
rect 15256 2148 15312 2150
rect 13266 584 13322 640
rect 12714 312 12770 368
rect 13542 448 13598 504
rect 14922 176 14978 232
rect 14646 40 14702 96
rect 15842 4256 15898 4312
rect 16854 3984 16910 4040
rect 15750 3304 15806 3360
rect 15566 1944 15622 2000
rect 17774 5228 17830 5264
rect 17774 5208 17776 5228
rect 17776 5208 17828 5228
rect 17828 5208 17830 5228
rect 17866 5072 17922 5128
rect 16302 1808 16358 1864
rect 16854 1672 16910 1728
rect 18602 3440 18658 3496
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 20196 6010 20252 6012
rect 19956 5958 20002 6010
rect 20002 5958 20012 6010
rect 20036 5958 20066 6010
rect 20066 5958 20078 6010
rect 20078 5958 20092 6010
rect 20116 5958 20130 6010
rect 20130 5958 20142 6010
rect 20142 5958 20172 6010
rect 20196 5958 20206 6010
rect 20206 5958 20252 6010
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 20196 5956 20252 5958
rect 21362 5772 21418 5808
rect 21362 5752 21364 5772
rect 21364 5752 21416 5772
rect 21416 5752 21418 5772
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 20196 4922 20252 4924
rect 19956 4870 20002 4922
rect 20002 4870 20012 4922
rect 20036 4870 20066 4922
rect 20066 4870 20078 4922
rect 20078 4870 20092 4922
rect 20116 4870 20130 4922
rect 20130 4870 20142 4922
rect 20142 4870 20172 4922
rect 20196 4870 20206 4922
rect 20206 4870 20252 4922
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 20196 4868 20252 4870
rect 19798 4256 19854 4312
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 20196 3834 20252 3836
rect 19956 3782 20002 3834
rect 20002 3782 20012 3834
rect 20036 3782 20066 3834
rect 20066 3782 20078 3834
rect 20078 3782 20092 3834
rect 20116 3782 20130 3834
rect 20130 3782 20142 3834
rect 20142 3782 20172 3834
rect 20196 3782 20206 3834
rect 20206 3782 20252 3834
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 20196 3780 20252 3782
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 20196 2746 20252 2748
rect 19956 2694 20002 2746
rect 20002 2694 20012 2746
rect 20036 2694 20066 2746
rect 20066 2694 20078 2746
rect 20078 2694 20092 2746
rect 20116 2694 20130 2746
rect 20130 2694 20142 2746
rect 20142 2694 20172 2746
rect 20196 2694 20206 2746
rect 20206 2694 20252 2746
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 20196 2692 20252 2694
rect 21016 5466 21072 5468
rect 21096 5466 21152 5468
rect 21176 5466 21232 5468
rect 21256 5466 21312 5468
rect 21016 5414 21062 5466
rect 21062 5414 21072 5466
rect 21096 5414 21126 5466
rect 21126 5414 21138 5466
rect 21138 5414 21152 5466
rect 21176 5414 21190 5466
rect 21190 5414 21202 5466
rect 21202 5414 21232 5466
rect 21256 5414 21266 5466
rect 21266 5414 21312 5466
rect 21016 5412 21072 5414
rect 21096 5412 21152 5414
rect 21176 5412 21232 5414
rect 21256 5412 21312 5414
rect 21362 4664 21418 4720
rect 21016 4378 21072 4380
rect 21096 4378 21152 4380
rect 21176 4378 21232 4380
rect 21256 4378 21312 4380
rect 21016 4326 21062 4378
rect 21062 4326 21072 4378
rect 21096 4326 21126 4378
rect 21126 4326 21138 4378
rect 21138 4326 21152 4378
rect 21176 4326 21190 4378
rect 21190 4326 21202 4378
rect 21202 4326 21232 4378
rect 21256 4326 21266 4378
rect 21266 4326 21312 4378
rect 21016 4324 21072 4326
rect 21096 4324 21152 4326
rect 21176 4324 21232 4326
rect 21256 4324 21312 4326
rect 20718 3984 20774 4040
rect 20534 1536 20590 1592
rect 21016 3290 21072 3292
rect 21096 3290 21152 3292
rect 21176 3290 21232 3292
rect 21256 3290 21312 3292
rect 21016 3238 21062 3290
rect 21062 3238 21072 3290
rect 21096 3238 21126 3290
rect 21126 3238 21138 3290
rect 21138 3238 21152 3290
rect 21176 3238 21190 3290
rect 21190 3238 21202 3290
rect 21202 3238 21232 3290
rect 21256 3238 21266 3290
rect 21266 3238 21312 3290
rect 21016 3236 21072 3238
rect 21096 3236 21152 3238
rect 21176 3236 21232 3238
rect 21256 3236 21312 3238
rect 20626 1128 20682 1184
rect 21016 2202 21072 2204
rect 21096 2202 21152 2204
rect 21176 2202 21232 2204
rect 21256 2202 21312 2204
rect 21016 2150 21062 2202
rect 21062 2150 21072 2202
rect 21096 2150 21126 2202
rect 21126 2150 21138 2202
rect 21138 2150 21152 2202
rect 21176 2150 21190 2202
rect 21190 2150 21202 2202
rect 21202 2150 21232 2202
rect 21256 2150 21266 2202
rect 21266 2150 21312 2202
rect 21016 2148 21072 2150
rect 21096 2148 21152 2150
rect 21176 2148 21232 2150
rect 21256 2148 21312 2150
rect 22282 6160 22338 6216
rect 22190 5616 22246 5672
rect 22006 4004 22062 4040
rect 22006 3984 22008 4004
rect 22008 3984 22060 4004
rect 22060 3984 22062 4004
rect 21822 3612 21824 3632
rect 21824 3612 21876 3632
rect 21876 3612 21878 3632
rect 21822 3576 21878 3612
rect 21730 2896 21786 2952
rect 22834 4528 22890 4584
rect 22558 1400 22614 1456
rect 23294 4120 23350 4176
rect 23018 3032 23074 3088
rect 23662 3732 23718 3768
rect 23662 3712 23664 3732
rect 23664 3712 23716 3732
rect 23716 3712 23718 3732
rect 23110 2760 23166 2816
rect 22926 2488 22982 2544
rect 24122 2488 24178 2544
rect 24214 584 24270 640
rect 24950 1672 25006 1728
rect 25042 312 25098 368
rect 25956 8186 26012 8188
rect 26036 8186 26092 8188
rect 26116 8186 26172 8188
rect 26196 8186 26252 8188
rect 25956 8134 26002 8186
rect 26002 8134 26012 8186
rect 26036 8134 26066 8186
rect 26066 8134 26078 8186
rect 26078 8134 26092 8186
rect 26116 8134 26130 8186
rect 26130 8134 26142 8186
rect 26142 8134 26172 8186
rect 26196 8134 26206 8186
rect 26206 8134 26252 8186
rect 25956 8132 26012 8134
rect 26036 8132 26092 8134
rect 26116 8132 26172 8134
rect 26196 8132 26252 8134
rect 26238 7384 26294 7440
rect 27016 8730 27072 8732
rect 27096 8730 27152 8732
rect 27176 8730 27232 8732
rect 27256 8730 27312 8732
rect 27016 8678 27062 8730
rect 27062 8678 27072 8730
rect 27096 8678 27126 8730
rect 27126 8678 27138 8730
rect 27138 8678 27152 8730
rect 27176 8678 27190 8730
rect 27190 8678 27202 8730
rect 27202 8678 27232 8730
rect 27256 8678 27266 8730
rect 27266 8678 27312 8730
rect 27016 8676 27072 8678
rect 27096 8676 27152 8678
rect 27176 8676 27232 8678
rect 27256 8676 27312 8678
rect 33016 8730 33072 8732
rect 33096 8730 33152 8732
rect 33176 8730 33232 8732
rect 33256 8730 33312 8732
rect 33016 8678 33062 8730
rect 33062 8678 33072 8730
rect 33096 8678 33126 8730
rect 33126 8678 33138 8730
rect 33138 8678 33152 8730
rect 33176 8678 33190 8730
rect 33190 8678 33202 8730
rect 33202 8678 33232 8730
rect 33256 8678 33266 8730
rect 33266 8678 33312 8730
rect 33016 8676 33072 8678
rect 33096 8676 33152 8678
rect 33176 8676 33232 8678
rect 33256 8676 33312 8678
rect 36358 9560 36414 9616
rect 36910 9288 36966 9344
rect 27016 7642 27072 7644
rect 27096 7642 27152 7644
rect 27176 7642 27232 7644
rect 27256 7642 27312 7644
rect 27016 7590 27062 7642
rect 27062 7590 27072 7642
rect 27096 7590 27126 7642
rect 27126 7590 27138 7642
rect 27138 7590 27152 7642
rect 27176 7590 27190 7642
rect 27190 7590 27202 7642
rect 27202 7590 27232 7642
rect 27256 7590 27266 7642
rect 27266 7590 27312 7642
rect 27016 7588 27072 7590
rect 27096 7588 27152 7590
rect 27176 7588 27232 7590
rect 27256 7588 27312 7590
rect 25956 7098 26012 7100
rect 26036 7098 26092 7100
rect 26116 7098 26172 7100
rect 26196 7098 26252 7100
rect 25956 7046 26002 7098
rect 26002 7046 26012 7098
rect 26036 7046 26066 7098
rect 26066 7046 26078 7098
rect 26078 7046 26092 7098
rect 26116 7046 26130 7098
rect 26130 7046 26142 7098
rect 26142 7046 26172 7098
rect 26196 7046 26206 7098
rect 26206 7046 26252 7098
rect 25956 7044 26012 7046
rect 26036 7044 26092 7046
rect 26116 7044 26172 7046
rect 26196 7044 26252 7046
rect 25956 6010 26012 6012
rect 26036 6010 26092 6012
rect 26116 6010 26172 6012
rect 26196 6010 26252 6012
rect 25956 5958 26002 6010
rect 26002 5958 26012 6010
rect 26036 5958 26066 6010
rect 26066 5958 26078 6010
rect 26078 5958 26092 6010
rect 26116 5958 26130 6010
rect 26130 5958 26142 6010
rect 26142 5958 26172 6010
rect 26196 5958 26206 6010
rect 26206 5958 26252 6010
rect 25956 5956 26012 5958
rect 26036 5956 26092 5958
rect 26116 5956 26172 5958
rect 26196 5956 26252 5958
rect 25956 4922 26012 4924
rect 26036 4922 26092 4924
rect 26116 4922 26172 4924
rect 26196 4922 26252 4924
rect 25956 4870 26002 4922
rect 26002 4870 26012 4922
rect 26036 4870 26066 4922
rect 26066 4870 26078 4922
rect 26078 4870 26092 4922
rect 26116 4870 26130 4922
rect 26130 4870 26142 4922
rect 26142 4870 26172 4922
rect 26196 4870 26206 4922
rect 26206 4870 26252 4922
rect 25956 4868 26012 4870
rect 26036 4868 26092 4870
rect 26116 4868 26172 4870
rect 26196 4868 26252 4870
rect 25956 3834 26012 3836
rect 26036 3834 26092 3836
rect 26116 3834 26172 3836
rect 26196 3834 26252 3836
rect 25956 3782 26002 3834
rect 26002 3782 26012 3834
rect 26036 3782 26066 3834
rect 26066 3782 26078 3834
rect 26078 3782 26092 3834
rect 26116 3782 26130 3834
rect 26130 3782 26142 3834
rect 26142 3782 26172 3834
rect 26196 3782 26206 3834
rect 26206 3782 26252 3834
rect 25956 3780 26012 3782
rect 26036 3780 26092 3782
rect 26116 3780 26172 3782
rect 26196 3780 26252 3782
rect 25956 2746 26012 2748
rect 26036 2746 26092 2748
rect 26116 2746 26172 2748
rect 26196 2746 26252 2748
rect 25956 2694 26002 2746
rect 26002 2694 26012 2746
rect 26036 2694 26066 2746
rect 26066 2694 26078 2746
rect 26078 2694 26092 2746
rect 26116 2694 26130 2746
rect 26130 2694 26142 2746
rect 26142 2694 26172 2746
rect 26196 2694 26206 2746
rect 26206 2694 26252 2746
rect 25956 2692 26012 2694
rect 26036 2692 26092 2694
rect 26116 2692 26172 2694
rect 26196 2692 26252 2694
rect 26146 448 26202 504
rect 27016 6554 27072 6556
rect 27096 6554 27152 6556
rect 27176 6554 27232 6556
rect 27256 6554 27312 6556
rect 27016 6502 27062 6554
rect 27062 6502 27072 6554
rect 27096 6502 27126 6554
rect 27126 6502 27138 6554
rect 27138 6502 27152 6554
rect 27176 6502 27190 6554
rect 27190 6502 27202 6554
rect 27202 6502 27232 6554
rect 27256 6502 27266 6554
rect 27266 6502 27312 6554
rect 27016 6500 27072 6502
rect 27096 6500 27152 6502
rect 27176 6500 27232 6502
rect 27256 6500 27312 6502
rect 27016 5466 27072 5468
rect 27096 5466 27152 5468
rect 27176 5466 27232 5468
rect 27256 5466 27312 5468
rect 27016 5414 27062 5466
rect 27062 5414 27072 5466
rect 27096 5414 27126 5466
rect 27126 5414 27138 5466
rect 27138 5414 27152 5466
rect 27176 5414 27190 5466
rect 27190 5414 27202 5466
rect 27202 5414 27232 5466
rect 27256 5414 27266 5466
rect 27266 5414 27312 5466
rect 27016 5412 27072 5414
rect 27096 5412 27152 5414
rect 27176 5412 27232 5414
rect 27256 5412 27312 5414
rect 27016 4378 27072 4380
rect 27096 4378 27152 4380
rect 27176 4378 27232 4380
rect 27256 4378 27312 4380
rect 27016 4326 27062 4378
rect 27062 4326 27072 4378
rect 27096 4326 27126 4378
rect 27126 4326 27138 4378
rect 27138 4326 27152 4378
rect 27176 4326 27190 4378
rect 27190 4326 27202 4378
rect 27202 4326 27232 4378
rect 27256 4326 27266 4378
rect 27266 4326 27312 4378
rect 27016 4324 27072 4326
rect 27096 4324 27152 4326
rect 27176 4324 27232 4326
rect 27256 4324 27312 4326
rect 27016 3290 27072 3292
rect 27096 3290 27152 3292
rect 27176 3290 27232 3292
rect 27256 3290 27312 3292
rect 27016 3238 27062 3290
rect 27062 3238 27072 3290
rect 27096 3238 27126 3290
rect 27126 3238 27138 3290
rect 27138 3238 27152 3290
rect 27176 3238 27190 3290
rect 27190 3238 27202 3290
rect 27202 3238 27232 3290
rect 27256 3238 27266 3290
rect 27266 3238 27312 3290
rect 27016 3236 27072 3238
rect 27096 3236 27152 3238
rect 27176 3236 27232 3238
rect 27256 3236 27312 3238
rect 27016 2202 27072 2204
rect 27096 2202 27152 2204
rect 27176 2202 27232 2204
rect 27256 2202 27312 2204
rect 27016 2150 27062 2202
rect 27062 2150 27072 2202
rect 27096 2150 27126 2202
rect 27126 2150 27138 2202
rect 27138 2150 27152 2202
rect 27176 2150 27190 2202
rect 27190 2150 27202 2202
rect 27202 2150 27232 2202
rect 27256 2150 27266 2202
rect 27266 2150 27312 2202
rect 27016 2148 27072 2150
rect 27096 2148 27152 2150
rect 27176 2148 27232 2150
rect 27256 2148 27312 2150
rect 28262 1808 28318 1864
rect 29274 3476 29276 3496
rect 29276 3476 29328 3496
rect 29328 3476 29330 3496
rect 29274 3440 29330 3476
rect 29366 176 29422 232
rect 29734 2352 29790 2408
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 33016 7642 33072 7644
rect 33096 7642 33152 7644
rect 33176 7642 33232 7644
rect 33256 7642 33312 7644
rect 33016 7590 33062 7642
rect 33062 7590 33072 7642
rect 33096 7590 33126 7642
rect 33126 7590 33138 7642
rect 33138 7590 33152 7642
rect 33176 7590 33190 7642
rect 33190 7590 33202 7642
rect 33202 7590 33232 7642
rect 33256 7590 33266 7642
rect 33266 7590 33312 7642
rect 33016 7588 33072 7590
rect 33096 7588 33152 7590
rect 33176 7588 33232 7590
rect 33256 7588 33312 7590
rect 31758 6160 31814 6216
rect 30838 40 30894 96
rect 31482 1400 31538 1456
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 33414 7384 33470 7440
rect 33016 6554 33072 6556
rect 33096 6554 33152 6556
rect 33176 6554 33232 6556
rect 33256 6554 33312 6556
rect 33016 6502 33062 6554
rect 33062 6502 33072 6554
rect 33096 6502 33126 6554
rect 33126 6502 33138 6554
rect 33138 6502 33152 6554
rect 33176 6502 33190 6554
rect 33190 6502 33202 6554
rect 33202 6502 33232 6554
rect 33256 6502 33266 6554
rect 33266 6502 33312 6554
rect 33016 6500 33072 6502
rect 33096 6500 33152 6502
rect 33176 6500 33232 6502
rect 33256 6500 33312 6502
rect 33016 5466 33072 5468
rect 33096 5466 33152 5468
rect 33176 5466 33232 5468
rect 33256 5466 33312 5468
rect 33016 5414 33062 5466
rect 33062 5414 33072 5466
rect 33096 5414 33126 5466
rect 33126 5414 33138 5466
rect 33138 5414 33152 5466
rect 33176 5414 33190 5466
rect 33190 5414 33202 5466
rect 33202 5414 33232 5466
rect 33256 5414 33266 5466
rect 33266 5414 33312 5466
rect 33016 5412 33072 5414
rect 33096 5412 33152 5414
rect 33176 5412 33232 5414
rect 33256 5412 33312 5414
rect 33016 4378 33072 4380
rect 33096 4378 33152 4380
rect 33176 4378 33232 4380
rect 33256 4378 33312 4380
rect 33016 4326 33062 4378
rect 33062 4326 33072 4378
rect 33096 4326 33126 4378
rect 33126 4326 33138 4378
rect 33138 4326 33152 4378
rect 33176 4326 33190 4378
rect 33190 4326 33202 4378
rect 33202 4326 33232 4378
rect 33256 4326 33266 4378
rect 33266 4326 33312 4378
rect 33016 4324 33072 4326
rect 33096 4324 33152 4326
rect 33176 4324 33232 4326
rect 33256 4324 33312 4326
rect 33016 3290 33072 3292
rect 33096 3290 33152 3292
rect 33176 3290 33232 3292
rect 33256 3290 33312 3292
rect 33016 3238 33062 3290
rect 33062 3238 33072 3290
rect 33096 3238 33126 3290
rect 33126 3238 33138 3290
rect 33138 3238 33152 3290
rect 33176 3238 33190 3290
rect 33190 3238 33202 3290
rect 33202 3238 33232 3290
rect 33256 3238 33266 3290
rect 33266 3238 33312 3290
rect 33016 3236 33072 3238
rect 33096 3236 33152 3238
rect 33176 3236 33232 3238
rect 33256 3236 33312 3238
rect 33138 2896 33194 2952
rect 32862 2488 32918 2544
rect 33016 2202 33072 2204
rect 33096 2202 33152 2204
rect 33176 2202 33232 2204
rect 33256 2202 33312 2204
rect 33016 2150 33062 2202
rect 33062 2150 33072 2202
rect 33096 2150 33126 2202
rect 33126 2150 33138 2202
rect 33138 2150 33152 2202
rect 33176 2150 33190 2202
rect 33190 2150 33202 2202
rect 33202 2150 33232 2202
rect 33256 2150 33266 2202
rect 33266 2150 33312 2202
rect 33016 2148 33072 2150
rect 33096 2148 33152 2150
rect 33176 2148 33232 2150
rect 33256 2148 33312 2150
rect 33506 3576 33562 3632
rect 37278 9016 37334 9072
rect 37646 8472 37702 8528
rect 38474 8744 38530 8800
rect 37956 8186 38012 8188
rect 38036 8186 38092 8188
rect 38116 8186 38172 8188
rect 38196 8186 38252 8188
rect 37956 8134 38002 8186
rect 38002 8134 38012 8186
rect 38036 8134 38066 8186
rect 38066 8134 38078 8186
rect 38078 8134 38092 8186
rect 38116 8134 38130 8186
rect 38130 8134 38142 8186
rect 38142 8134 38172 8186
rect 38196 8134 38206 8186
rect 38206 8134 38252 8186
rect 37956 8132 38012 8134
rect 38036 8132 38092 8134
rect 38116 8132 38172 8134
rect 38196 8132 38252 8134
rect 38382 7692 38384 7712
rect 38384 7692 38436 7712
rect 38436 7692 38438 7712
rect 38382 7656 38438 7692
rect 38750 8200 38806 8256
rect 38934 7928 38990 7984
rect 38014 7384 38070 7440
rect 38382 7148 38384 7168
rect 38384 7148 38436 7168
rect 38436 7148 38438 7168
rect 38382 7112 38438 7148
rect 37956 7098 38012 7100
rect 38036 7098 38092 7100
rect 38116 7098 38172 7100
rect 38196 7098 38252 7100
rect 37956 7046 38002 7098
rect 38002 7046 38012 7098
rect 38036 7046 38066 7098
rect 38066 7046 38078 7098
rect 38078 7046 38092 7098
rect 38116 7046 38130 7098
rect 38130 7046 38142 7098
rect 38142 7046 38172 7098
rect 38196 7046 38206 7098
rect 38206 7046 38252 7098
rect 37956 7044 38012 7046
rect 38036 7044 38092 7046
rect 38116 7044 38172 7046
rect 38196 7044 38252 7046
rect 38198 6840 38254 6896
rect 38382 6840 38438 6896
rect 38014 6604 38016 6624
rect 38016 6604 38068 6624
rect 38068 6604 38070 6624
rect 38014 6568 38070 6604
rect 38382 6296 38438 6352
rect 35898 3984 35954 4040
rect 39118 6060 39120 6080
rect 39120 6060 39172 6080
rect 39172 6060 39174 6080
rect 39118 6024 39174 6060
rect 37956 6010 38012 6012
rect 38036 6010 38092 6012
rect 38116 6010 38172 6012
rect 38196 6010 38252 6012
rect 37956 5958 38002 6010
rect 38002 5958 38012 6010
rect 38036 5958 38066 6010
rect 38066 5958 38078 6010
rect 38078 5958 38092 6010
rect 38116 5958 38130 6010
rect 38130 5958 38142 6010
rect 38142 5958 38172 6010
rect 38196 5958 38206 6010
rect 38206 5958 38252 6010
rect 37956 5956 38012 5958
rect 38036 5956 38092 5958
rect 38116 5956 38172 5958
rect 38196 5956 38252 5958
rect 38382 5788 38384 5808
rect 38384 5788 38436 5808
rect 38436 5788 38438 5808
rect 38382 5752 38438 5788
rect 36634 1944 36690 2000
rect 38014 5516 38016 5536
rect 38016 5516 38068 5536
rect 38068 5516 38070 5536
rect 38014 5480 38070 5516
rect 38382 5208 38438 5264
rect 39118 4972 39120 4992
rect 39120 4972 39172 4992
rect 39172 4972 39174 4992
rect 39118 4936 39174 4972
rect 37956 4922 38012 4924
rect 38036 4922 38092 4924
rect 38116 4922 38172 4924
rect 38196 4922 38252 4924
rect 37956 4870 38002 4922
rect 38002 4870 38012 4922
rect 38036 4870 38066 4922
rect 38066 4870 38078 4922
rect 38078 4870 38092 4922
rect 38116 4870 38130 4922
rect 38130 4870 38142 4922
rect 38142 4870 38172 4922
rect 38196 4870 38206 4922
rect 38206 4870 38252 4922
rect 37956 4868 38012 4870
rect 38036 4868 38092 4870
rect 38116 4868 38172 4870
rect 38196 4868 38252 4870
rect 38382 4700 38384 4720
rect 38384 4700 38436 4720
rect 38436 4700 38438 4720
rect 38014 4428 38016 4448
rect 38016 4428 38068 4448
rect 38068 4428 38070 4448
rect 38014 4392 38070 4428
rect 38382 4664 38438 4700
rect 38382 4120 38438 4176
rect 39118 3884 39120 3904
rect 39120 3884 39172 3904
rect 39172 3884 39174 3904
rect 39118 3848 39174 3884
rect 37956 3834 38012 3836
rect 38036 3834 38092 3836
rect 38116 3834 38172 3836
rect 38196 3834 38252 3836
rect 37956 3782 38002 3834
rect 38002 3782 38012 3834
rect 38036 3782 38066 3834
rect 38066 3782 38078 3834
rect 38078 3782 38092 3834
rect 38116 3782 38130 3834
rect 38130 3782 38142 3834
rect 38142 3782 38172 3834
rect 38196 3782 38206 3834
rect 38206 3782 38252 3834
rect 37956 3780 38012 3782
rect 38036 3780 38092 3782
rect 38116 3780 38172 3782
rect 38196 3780 38252 3782
rect 38382 3612 38384 3632
rect 38384 3612 38436 3632
rect 38436 3612 38438 3632
rect 38382 3576 38438 3612
rect 38014 3340 38016 3360
rect 38016 3340 38068 3360
rect 38068 3340 38070 3360
rect 38014 3304 38070 3340
rect 38382 3032 38438 3088
rect 39118 2796 39120 2816
rect 39120 2796 39172 2816
rect 39172 2796 39174 2816
rect 37186 1400 37242 1456
rect 39118 2760 39174 2796
rect 37956 2746 38012 2748
rect 38036 2746 38092 2748
rect 38116 2746 38172 2748
rect 38196 2746 38252 2748
rect 37956 2694 38002 2746
rect 38002 2694 38012 2746
rect 38036 2694 38066 2746
rect 38066 2694 38078 2746
rect 38078 2694 38092 2746
rect 38116 2694 38130 2746
rect 38130 2694 38142 2746
rect 38142 2694 38172 2746
rect 38196 2694 38206 2746
rect 38206 2694 38252 2746
rect 37956 2692 38012 2694
rect 38036 2692 38092 2694
rect 38116 2692 38172 2694
rect 38196 2692 38252 2694
rect 38382 2524 38384 2544
rect 38384 2524 38436 2544
rect 38436 2524 38438 2544
rect 38382 2488 38438 2524
rect 38014 2252 38016 2272
rect 38016 2252 38068 2272
rect 38068 2252 38070 2272
rect 38014 2216 38070 2252
rect 37830 1672 37886 1728
rect 37646 1128 37702 1184
<< metal3 >>
rect 0 9618 120 9648
rect 19793 9618 19859 9621
rect 0 9616 19859 9618
rect 0 9560 19798 9616
rect 19854 9560 19859 9616
rect 0 9558 19859 9560
rect 0 9528 120 9558
rect 19793 9555 19859 9558
rect 36353 9618 36419 9621
rect 39808 9618 39928 9648
rect 36353 9616 39928 9618
rect 36353 9560 36358 9616
rect 36414 9560 39928 9616
rect 36353 9558 39928 9560
rect 36353 9555 36419 9558
rect 39808 9528 39928 9558
rect 0 9346 120 9376
rect 14641 9346 14707 9349
rect 0 9344 14707 9346
rect 0 9288 14646 9344
rect 14702 9288 14707 9344
rect 0 9286 14707 9288
rect 0 9256 120 9286
rect 14641 9283 14707 9286
rect 36905 9346 36971 9349
rect 39808 9346 39928 9376
rect 36905 9344 39928 9346
rect 36905 9288 36910 9344
rect 36966 9288 39928 9344
rect 36905 9286 39928 9288
rect 36905 9283 36971 9286
rect 39808 9256 39928 9286
rect 0 9074 120 9104
rect 14825 9074 14891 9077
rect 0 9072 14891 9074
rect 0 9016 14830 9072
rect 14886 9016 14891 9072
rect 0 9014 14891 9016
rect 0 8984 120 9014
rect 14825 9011 14891 9014
rect 37273 9074 37339 9077
rect 39808 9074 39928 9104
rect 37273 9072 39928 9074
rect 37273 9016 37278 9072
rect 37334 9016 39928 9072
rect 37273 9014 39928 9016
rect 37273 9011 37339 9014
rect 39808 8984 39928 9014
rect 0 8802 120 8832
rect 2865 8802 2931 8805
rect 0 8800 2931 8802
rect 0 8744 2870 8800
rect 2926 8744 2931 8800
rect 0 8742 2931 8744
rect 0 8712 120 8742
rect 2865 8739 2931 8742
rect 38469 8802 38535 8805
rect 39808 8802 39928 8832
rect 38469 8800 39928 8802
rect 38469 8744 38474 8800
rect 38530 8744 39928 8800
rect 38469 8742 39928 8744
rect 38469 8739 38535 8742
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 9006 8736 9322 8737
rect 9006 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9322 8736
rect 9006 8671 9322 8672
rect 15006 8736 15322 8737
rect 15006 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15322 8736
rect 15006 8671 15322 8672
rect 21006 8736 21322 8737
rect 21006 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21322 8736
rect 21006 8671 21322 8672
rect 27006 8736 27322 8737
rect 27006 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27322 8736
rect 27006 8671 27322 8672
rect 33006 8736 33322 8737
rect 33006 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33322 8736
rect 39808 8712 39928 8742
rect 33006 8671 33322 8672
rect 0 8530 120 8560
rect 17033 8530 17099 8533
rect 0 8528 17099 8530
rect 0 8472 17038 8528
rect 17094 8472 17099 8528
rect 0 8470 17099 8472
rect 0 8440 120 8470
rect 17033 8467 17099 8470
rect 37641 8530 37707 8533
rect 39808 8530 39928 8560
rect 37641 8528 39928 8530
rect 37641 8472 37646 8528
rect 37702 8472 39928 8528
rect 37641 8470 39928 8472
rect 37641 8467 37707 8470
rect 39808 8440 39928 8470
rect 2865 8394 2931 8397
rect 14917 8394 14983 8397
rect 2865 8392 14983 8394
rect 2865 8336 2870 8392
rect 2926 8336 14922 8392
rect 14978 8336 14983 8392
rect 2865 8334 14983 8336
rect 2865 8331 2931 8334
rect 14917 8331 14983 8334
rect 0 8258 120 8288
rect 1761 8258 1827 8261
rect 0 8256 1827 8258
rect 0 8200 1766 8256
rect 1822 8200 1827 8256
rect 0 8198 1827 8200
rect 0 8168 120 8198
rect 1761 8195 1827 8198
rect 38745 8258 38811 8261
rect 39808 8258 39928 8288
rect 38745 8256 39928 8258
rect 38745 8200 38750 8256
rect 38806 8200 39928 8256
rect 38745 8198 39928 8200
rect 38745 8195 38811 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 7946 8127 8262 8128
rect 13946 8192 14262 8193
rect 13946 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14262 8192
rect 13946 8127 14262 8128
rect 19946 8192 20262 8193
rect 19946 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20262 8192
rect 19946 8127 20262 8128
rect 25946 8192 26262 8193
rect 25946 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26262 8192
rect 25946 8127 26262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 31946 8127 32262 8128
rect 37946 8192 38262 8193
rect 37946 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38262 8192
rect 39808 8168 39928 8198
rect 37946 8127 38262 8128
rect 0 7986 120 8016
rect 18229 7986 18295 7989
rect 0 7984 18295 7986
rect 0 7928 18234 7984
rect 18290 7928 18295 7984
rect 0 7926 18295 7928
rect 0 7896 120 7926
rect 18229 7923 18295 7926
rect 38929 7986 38995 7989
rect 39808 7986 39928 8016
rect 38929 7984 39928 7986
rect 38929 7928 38934 7984
rect 38990 7928 39928 7984
rect 38929 7926 39928 7928
rect 38929 7923 38995 7926
rect 39808 7896 39928 7926
rect 18045 7850 18111 7853
rect 18597 7850 18663 7853
rect 2730 7848 18663 7850
rect 2730 7792 18050 7848
rect 18106 7792 18602 7848
rect 18658 7792 18663 7848
rect 2730 7790 18663 7792
rect 0 7714 120 7744
rect 2730 7714 2790 7790
rect 18045 7787 18111 7790
rect 18597 7787 18663 7790
rect 0 7654 2790 7714
rect 38377 7714 38443 7717
rect 39808 7714 39928 7744
rect 38377 7712 39928 7714
rect 38377 7656 38382 7712
rect 38438 7656 39928 7712
rect 38377 7654 39928 7656
rect 0 7624 120 7654
rect 38377 7651 38443 7654
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 9006 7648 9322 7649
rect 9006 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9322 7648
rect 9006 7583 9322 7584
rect 15006 7648 15322 7649
rect 15006 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15322 7648
rect 15006 7583 15322 7584
rect 21006 7648 21322 7649
rect 21006 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21322 7648
rect 21006 7583 21322 7584
rect 27006 7648 27322 7649
rect 27006 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27322 7648
rect 27006 7583 27322 7584
rect 33006 7648 33322 7649
rect 33006 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33322 7648
rect 39808 7624 39928 7654
rect 33006 7583 33322 7584
rect 0 7442 120 7472
rect 15285 7442 15351 7445
rect 0 7440 15351 7442
rect 0 7384 15290 7440
rect 15346 7384 15351 7440
rect 0 7382 15351 7384
rect 0 7352 120 7382
rect 15285 7379 15351 7382
rect 26233 7442 26299 7445
rect 33409 7442 33475 7445
rect 26233 7440 33475 7442
rect 26233 7384 26238 7440
rect 26294 7384 33414 7440
rect 33470 7384 33475 7440
rect 26233 7382 33475 7384
rect 26233 7379 26299 7382
rect 33409 7379 33475 7382
rect 38009 7442 38075 7445
rect 39808 7442 39928 7472
rect 38009 7440 39928 7442
rect 38009 7384 38014 7440
rect 38070 7384 39928 7440
rect 38009 7382 39928 7384
rect 38009 7379 38075 7382
rect 39808 7352 39928 7382
rect 1761 7306 1827 7309
rect 19517 7306 19583 7309
rect 20253 7306 20319 7309
rect 1761 7304 20319 7306
rect 1761 7248 1766 7304
rect 1822 7248 19522 7304
rect 19578 7248 20258 7304
rect 20314 7248 20319 7304
rect 1761 7246 20319 7248
rect 1761 7243 1827 7246
rect 19517 7243 19583 7246
rect 20253 7243 20319 7246
rect 0 7170 120 7200
rect 1301 7170 1367 7173
rect 0 7168 1367 7170
rect 0 7112 1306 7168
rect 1362 7112 1367 7168
rect 0 7110 1367 7112
rect 0 7080 120 7110
rect 1301 7107 1367 7110
rect 38377 7170 38443 7173
rect 39808 7170 39928 7200
rect 38377 7168 39928 7170
rect 38377 7112 38382 7168
rect 38438 7112 39928 7168
rect 38377 7110 39928 7112
rect 38377 7107 38443 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 7946 7039 8262 7040
rect 13946 7104 14262 7105
rect 13946 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14262 7104
rect 13946 7039 14262 7040
rect 19946 7104 20262 7105
rect 19946 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20262 7104
rect 19946 7039 20262 7040
rect 25946 7104 26262 7105
rect 25946 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26262 7104
rect 25946 7039 26262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 31946 7039 32262 7040
rect 37946 7104 38262 7105
rect 37946 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38262 7104
rect 39808 7080 39928 7110
rect 37946 7039 38262 7040
rect 0 6898 120 6928
rect 15745 6898 15811 6901
rect 0 6896 15811 6898
rect 0 6840 15750 6896
rect 15806 6840 15811 6896
rect 0 6838 15811 6840
rect 0 6808 120 6838
rect 15745 6835 15811 6838
rect 16113 6898 16179 6901
rect 38193 6898 38259 6901
rect 16113 6896 38259 6898
rect 16113 6840 16118 6896
rect 16174 6840 38198 6896
rect 38254 6840 38259 6896
rect 16113 6838 38259 6840
rect 16113 6835 16179 6838
rect 38193 6835 38259 6838
rect 38377 6898 38443 6901
rect 39808 6898 39928 6928
rect 38377 6896 39928 6898
rect 38377 6840 38382 6896
rect 38438 6840 39928 6896
rect 38377 6838 39928 6840
rect 38377 6835 38443 6838
rect 39808 6808 39928 6838
rect 16665 6762 16731 6765
rect 2730 6760 16731 6762
rect 2730 6704 16670 6760
rect 16726 6704 16731 6760
rect 2730 6702 16731 6704
rect 0 6626 120 6656
rect 2730 6626 2790 6702
rect 16665 6699 16731 6702
rect 0 6566 2790 6626
rect 38009 6626 38075 6629
rect 39808 6626 39928 6656
rect 38009 6624 39928 6626
rect 38009 6568 38014 6624
rect 38070 6568 39928 6624
rect 38009 6566 39928 6568
rect 0 6536 120 6566
rect 38009 6563 38075 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 9006 6560 9322 6561
rect 9006 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9322 6560
rect 9006 6495 9322 6496
rect 15006 6560 15322 6561
rect 15006 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15322 6560
rect 15006 6495 15322 6496
rect 21006 6560 21322 6561
rect 21006 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21322 6560
rect 21006 6495 21322 6496
rect 27006 6560 27322 6561
rect 27006 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27322 6560
rect 27006 6495 27322 6496
rect 33006 6560 33322 6561
rect 33006 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33322 6560
rect 39808 6536 39928 6566
rect 33006 6495 33322 6496
rect 0 6354 120 6384
rect 18689 6354 18755 6357
rect 0 6352 18755 6354
rect 0 6296 18694 6352
rect 18750 6296 18755 6352
rect 0 6294 18755 6296
rect 0 6264 120 6294
rect 18689 6291 18755 6294
rect 38377 6354 38443 6357
rect 39808 6354 39928 6384
rect 38377 6352 39928 6354
rect 38377 6296 38382 6352
rect 38438 6296 39928 6352
rect 38377 6294 39928 6296
rect 38377 6291 38443 6294
rect 39808 6264 39928 6294
rect 17401 6218 17467 6221
rect 1764 6216 17467 6218
rect 1764 6160 17406 6216
rect 17462 6160 17467 6216
rect 1764 6158 17467 6160
rect 0 6082 120 6112
rect 1764 6082 1824 6158
rect 17401 6155 17467 6158
rect 22277 6218 22343 6221
rect 31753 6218 31819 6221
rect 22277 6216 31819 6218
rect 22277 6160 22282 6216
rect 22338 6160 31758 6216
rect 31814 6160 31819 6216
rect 22277 6158 31819 6160
rect 22277 6155 22343 6158
rect 31753 6155 31819 6158
rect 0 6022 1824 6082
rect 39113 6082 39179 6085
rect 39808 6082 39928 6112
rect 39113 6080 39928 6082
rect 39113 6024 39118 6080
rect 39174 6024 39928 6080
rect 39113 6022 39928 6024
rect 0 5992 120 6022
rect 39113 6019 39179 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 7946 5951 8262 5952
rect 13946 6016 14262 6017
rect 13946 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14262 6016
rect 13946 5951 14262 5952
rect 19946 6016 20262 6017
rect 19946 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20262 6016
rect 19946 5951 20262 5952
rect 25946 6016 26262 6017
rect 25946 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26262 6016
rect 25946 5951 26262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 31946 5951 32262 5952
rect 37946 6016 38262 6017
rect 37946 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38262 6016
rect 39808 5992 39928 6022
rect 37946 5951 38262 5952
rect 0 5810 120 5840
rect 21357 5810 21423 5813
rect 0 5808 21423 5810
rect 0 5752 21362 5808
rect 21418 5752 21423 5808
rect 0 5750 21423 5752
rect 0 5720 120 5750
rect 21357 5747 21423 5750
rect 38377 5810 38443 5813
rect 39808 5810 39928 5840
rect 38377 5808 39928 5810
rect 38377 5752 38382 5808
rect 38438 5752 39928 5808
rect 38377 5750 39928 5752
rect 38377 5747 38443 5750
rect 39808 5720 39928 5750
rect 3877 5674 3943 5677
rect 8293 5674 8359 5677
rect 3877 5672 8359 5674
rect 3877 5616 3882 5672
rect 3938 5616 8298 5672
rect 8354 5616 8359 5672
rect 3877 5614 8359 5616
rect 3877 5611 3943 5614
rect 8293 5611 8359 5614
rect 9949 5674 10015 5677
rect 22185 5674 22251 5677
rect 9949 5672 22251 5674
rect 9949 5616 9954 5672
rect 10010 5616 22190 5672
rect 22246 5616 22251 5672
rect 9949 5614 22251 5616
rect 9949 5611 10015 5614
rect 22185 5611 22251 5614
rect 0 5538 120 5568
rect 2865 5538 2931 5541
rect 0 5536 2931 5538
rect 0 5480 2870 5536
rect 2926 5480 2931 5536
rect 0 5478 2931 5480
rect 0 5448 120 5478
rect 2865 5475 2931 5478
rect 38009 5538 38075 5541
rect 39808 5538 39928 5568
rect 38009 5536 39928 5538
rect 38009 5480 38014 5536
rect 38070 5480 39928 5536
rect 38009 5478 39928 5480
rect 38009 5475 38075 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 9006 5472 9322 5473
rect 9006 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9322 5472
rect 9006 5407 9322 5408
rect 15006 5472 15322 5473
rect 15006 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15322 5472
rect 15006 5407 15322 5408
rect 21006 5472 21322 5473
rect 21006 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21322 5472
rect 21006 5407 21322 5408
rect 27006 5472 27322 5473
rect 27006 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27322 5472
rect 27006 5407 27322 5408
rect 33006 5472 33322 5473
rect 33006 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33322 5472
rect 39808 5448 39928 5478
rect 33006 5407 33322 5408
rect 0 5266 120 5296
rect 2773 5266 2839 5269
rect 0 5264 2839 5266
rect 0 5208 2778 5264
rect 2834 5208 2839 5264
rect 0 5206 2839 5208
rect 0 5176 120 5206
rect 2773 5203 2839 5206
rect 2957 5266 3023 5269
rect 17769 5266 17835 5269
rect 2957 5264 17835 5266
rect 2957 5208 2962 5264
rect 3018 5208 17774 5264
rect 17830 5208 17835 5264
rect 2957 5206 17835 5208
rect 2957 5203 3023 5206
rect 17769 5203 17835 5206
rect 38377 5266 38443 5269
rect 39808 5266 39928 5296
rect 38377 5264 39928 5266
rect 38377 5208 38382 5264
rect 38438 5208 39928 5264
rect 38377 5206 39928 5208
rect 38377 5203 38443 5206
rect 39808 5176 39928 5206
rect 2957 5130 3023 5133
rect 17861 5130 17927 5133
rect 1764 5070 2882 5130
rect 0 4994 120 5024
rect 1764 4994 1824 5070
rect 0 4934 1824 4994
rect 2822 4994 2882 5070
rect 2957 5128 17927 5130
rect 2957 5072 2962 5128
rect 3018 5072 17866 5128
rect 17922 5072 17927 5128
rect 2957 5070 17927 5072
rect 2957 5067 3023 5070
rect 17861 5067 17927 5070
rect 7649 4994 7715 4997
rect 2822 4992 7715 4994
rect 2822 4936 7654 4992
rect 7710 4936 7715 4992
rect 2822 4934 7715 4936
rect 0 4904 120 4934
rect 7649 4931 7715 4934
rect 39113 4994 39179 4997
rect 39808 4994 39928 5024
rect 39113 4992 39928 4994
rect 39113 4936 39118 4992
rect 39174 4936 39928 4992
rect 39113 4934 39928 4936
rect 39113 4931 39179 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 13946 4928 14262 4929
rect 13946 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14262 4928
rect 13946 4863 14262 4864
rect 19946 4928 20262 4929
rect 19946 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20262 4928
rect 19946 4863 20262 4864
rect 25946 4928 26262 4929
rect 25946 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26262 4928
rect 25946 4863 26262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 31946 4863 32262 4864
rect 37946 4928 38262 4929
rect 37946 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38262 4928
rect 39808 4904 39928 4934
rect 37946 4863 38262 4864
rect 0 4722 120 4752
rect 21357 4722 21423 4725
rect 0 4720 21423 4722
rect 0 4664 21362 4720
rect 21418 4664 21423 4720
rect 0 4662 21423 4664
rect 0 4632 120 4662
rect 21357 4659 21423 4662
rect 38377 4722 38443 4725
rect 39808 4722 39928 4752
rect 38377 4720 39928 4722
rect 38377 4664 38382 4720
rect 38438 4664 39928 4720
rect 38377 4662 39928 4664
rect 38377 4659 38443 4662
rect 39808 4632 39928 4662
rect 22829 4586 22895 4589
rect 2730 4584 22895 4586
rect 2730 4528 22834 4584
rect 22890 4528 22895 4584
rect 2730 4526 22895 4528
rect 0 4450 120 4480
rect 2730 4450 2790 4526
rect 22829 4523 22895 4526
rect 0 4390 2790 4450
rect 4429 4450 4495 4453
rect 8385 4450 8451 4453
rect 4429 4448 8451 4450
rect 4429 4392 4434 4448
rect 4490 4392 8390 4448
rect 8446 4392 8451 4448
rect 4429 4390 8451 4392
rect 0 4360 120 4390
rect 4429 4387 4495 4390
rect 8385 4387 8451 4390
rect 38009 4450 38075 4453
rect 39808 4450 39928 4480
rect 38009 4448 39928 4450
rect 38009 4392 38014 4448
rect 38070 4392 39928 4448
rect 38009 4390 39928 4392
rect 38009 4387 38075 4390
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 9006 4384 9322 4385
rect 9006 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9322 4384
rect 9006 4319 9322 4320
rect 15006 4384 15322 4385
rect 15006 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15322 4384
rect 15006 4319 15322 4320
rect 21006 4384 21322 4385
rect 21006 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21322 4384
rect 21006 4319 21322 4320
rect 27006 4384 27322 4385
rect 27006 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27322 4384
rect 27006 4319 27322 4320
rect 33006 4384 33322 4385
rect 33006 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33322 4384
rect 39808 4360 39928 4390
rect 33006 4319 33322 4320
rect 15837 4314 15903 4317
rect 19793 4314 19859 4317
rect 15837 4312 19859 4314
rect 15837 4256 15842 4312
rect 15898 4256 19798 4312
rect 19854 4256 19859 4312
rect 15837 4254 19859 4256
rect 15837 4251 15903 4254
rect 19793 4251 19859 4254
rect 0 4178 120 4208
rect 23289 4178 23355 4181
rect 0 4176 23355 4178
rect 0 4120 23294 4176
rect 23350 4120 23355 4176
rect 0 4118 23355 4120
rect 0 4088 120 4118
rect 23289 4115 23355 4118
rect 38377 4178 38443 4181
rect 39808 4178 39928 4208
rect 38377 4176 39928 4178
rect 38377 4120 38382 4176
rect 38438 4120 39928 4176
rect 38377 4118 39928 4120
rect 38377 4115 38443 4118
rect 39808 4088 39928 4118
rect 11053 4042 11119 4045
rect 16849 4042 16915 4045
rect 20713 4042 20779 4045
rect 1764 4040 11119 4042
rect 1764 3984 11058 4040
rect 11114 3984 11119 4040
rect 1764 3982 11119 3984
rect 0 3906 120 3936
rect 1764 3906 1824 3982
rect 11053 3979 11119 3982
rect 12390 4040 16915 4042
rect 12390 3984 16854 4040
rect 16910 3984 16915 4040
rect 12390 3982 16915 3984
rect 0 3846 1824 3906
rect 8753 3906 8819 3909
rect 12390 3906 12450 3982
rect 16849 3979 16915 3982
rect 19750 4040 20779 4042
rect 19750 3984 20718 4040
rect 20774 3984 20779 4040
rect 19750 3982 20779 3984
rect 19750 3906 19810 3982
rect 20713 3979 20779 3982
rect 22001 4042 22067 4045
rect 35893 4042 35959 4045
rect 22001 4040 35959 4042
rect 22001 3984 22006 4040
rect 22062 3984 35898 4040
rect 35954 3984 35959 4040
rect 22001 3982 35959 3984
rect 22001 3979 22067 3982
rect 35893 3979 35959 3982
rect 8753 3904 12450 3906
rect 8753 3848 8758 3904
rect 8814 3848 12450 3904
rect 8753 3846 12450 3848
rect 14414 3846 19810 3906
rect 39113 3906 39179 3909
rect 39808 3906 39928 3936
rect 39113 3904 39928 3906
rect 39113 3848 39118 3904
rect 39174 3848 39928 3904
rect 39113 3846 39928 3848
rect 0 3816 120 3846
rect 8753 3843 8819 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 13946 3840 14262 3841
rect 13946 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14262 3840
rect 13946 3775 14262 3776
rect 0 3634 120 3664
rect 14414 3634 14474 3846
rect 39113 3843 39179 3846
rect 19946 3840 20262 3841
rect 19946 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20262 3840
rect 19946 3775 20262 3776
rect 25946 3840 26262 3841
rect 25946 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26262 3840
rect 25946 3775 26262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 31946 3775 32262 3776
rect 37946 3840 38262 3841
rect 37946 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38262 3840
rect 39808 3816 39928 3846
rect 37946 3775 38262 3776
rect 23657 3770 23723 3773
rect 20486 3768 23723 3770
rect 20486 3712 23662 3768
rect 23718 3712 23723 3768
rect 20486 3710 23723 3712
rect 20486 3634 20546 3710
rect 23657 3707 23723 3710
rect 0 3574 14474 3634
rect 14598 3574 20546 3634
rect 21817 3634 21883 3637
rect 33501 3634 33567 3637
rect 21817 3632 33567 3634
rect 21817 3576 21822 3632
rect 21878 3576 33506 3632
rect 33562 3576 33567 3632
rect 21817 3574 33567 3576
rect 0 3544 120 3574
rect 14598 3498 14658 3574
rect 21817 3571 21883 3574
rect 33501 3571 33567 3574
rect 38377 3634 38443 3637
rect 39808 3634 39928 3664
rect 38377 3632 39928 3634
rect 38377 3576 38382 3632
rect 38438 3576 39928 3632
rect 38377 3574 39928 3576
rect 38377 3571 38443 3574
rect 39808 3544 39928 3574
rect 18597 3498 18663 3501
rect 29269 3498 29335 3501
rect 2730 3438 14658 3498
rect 14782 3496 18663 3498
rect 14782 3440 18602 3496
rect 18658 3440 18663 3496
rect 14782 3438 18663 3440
rect 0 3362 120 3392
rect 2730 3362 2790 3438
rect 0 3302 2790 3362
rect 0 3272 120 3302
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 9006 3296 9322 3297
rect 9006 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9322 3296
rect 9006 3231 9322 3232
rect 11145 3226 11211 3229
rect 14782 3226 14842 3438
rect 18597 3435 18663 3438
rect 18830 3496 29335 3498
rect 18830 3440 29274 3496
rect 29330 3440 29335 3496
rect 18830 3438 29335 3440
rect 15745 3362 15811 3365
rect 18830 3362 18890 3438
rect 29269 3435 29335 3438
rect 15745 3360 18890 3362
rect 15745 3304 15750 3360
rect 15806 3304 18890 3360
rect 15745 3302 18890 3304
rect 38009 3362 38075 3365
rect 39808 3362 39928 3392
rect 38009 3360 39928 3362
rect 38009 3304 38014 3360
rect 38070 3304 39928 3360
rect 38009 3302 39928 3304
rect 15745 3299 15811 3302
rect 38009 3299 38075 3302
rect 15006 3296 15322 3297
rect 15006 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15322 3296
rect 15006 3231 15322 3232
rect 21006 3296 21322 3297
rect 21006 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21322 3296
rect 21006 3231 21322 3232
rect 27006 3296 27322 3297
rect 27006 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27322 3296
rect 27006 3231 27322 3232
rect 33006 3296 33322 3297
rect 33006 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33322 3296
rect 39808 3272 39928 3302
rect 33006 3231 33322 3232
rect 11145 3224 14842 3226
rect 11145 3168 11150 3224
rect 11206 3168 14842 3224
rect 11145 3166 14842 3168
rect 11145 3163 11211 3166
rect 0 3090 120 3120
rect 23013 3090 23079 3093
rect 0 3088 23079 3090
rect 0 3032 23018 3088
rect 23074 3032 23079 3088
rect 0 3030 23079 3032
rect 0 3000 120 3030
rect 23013 3027 23079 3030
rect 38377 3090 38443 3093
rect 39808 3090 39928 3120
rect 38377 3088 39928 3090
rect 38377 3032 38382 3088
rect 38438 3032 39928 3088
rect 38377 3030 39928 3032
rect 38377 3027 38443 3030
rect 39808 3000 39928 3030
rect 21725 2954 21791 2957
rect 33133 2954 33199 2957
rect 1764 2894 20546 2954
rect 0 2818 120 2848
rect 1764 2818 1824 2894
rect 0 2758 1824 2818
rect 20486 2818 20546 2894
rect 21725 2952 33199 2954
rect 21725 2896 21730 2952
rect 21786 2896 33138 2952
rect 33194 2896 33199 2952
rect 21725 2894 33199 2896
rect 21725 2891 21791 2894
rect 33133 2891 33199 2894
rect 23105 2818 23171 2821
rect 20486 2816 23171 2818
rect 20486 2760 23110 2816
rect 23166 2760 23171 2816
rect 20486 2758 23171 2760
rect 0 2728 120 2758
rect 23105 2755 23171 2758
rect 39113 2818 39179 2821
rect 39808 2818 39928 2848
rect 39113 2816 39928 2818
rect 39113 2760 39118 2816
rect 39174 2760 39928 2816
rect 39113 2758 39928 2760
rect 39113 2755 39179 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 13946 2752 14262 2753
rect 13946 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14262 2752
rect 13946 2687 14262 2688
rect 19946 2752 20262 2753
rect 19946 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20262 2752
rect 19946 2687 20262 2688
rect 25946 2752 26262 2753
rect 25946 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26262 2752
rect 25946 2687 26262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 31946 2687 32262 2688
rect 37946 2752 38262 2753
rect 37946 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38262 2752
rect 39808 2728 39928 2758
rect 37946 2687 38262 2688
rect 11605 2682 11671 2685
rect 13169 2682 13235 2685
rect 11605 2680 13235 2682
rect 11605 2624 11610 2680
rect 11666 2624 13174 2680
rect 13230 2624 13235 2680
rect 11605 2622 13235 2624
rect 11605 2619 11671 2622
rect 13169 2619 13235 2622
rect 0 2546 120 2576
rect 565 2546 631 2549
rect 0 2544 631 2546
rect 0 2488 570 2544
rect 626 2488 631 2544
rect 0 2486 631 2488
rect 0 2456 120 2486
rect 565 2483 631 2486
rect 11881 2546 11947 2549
rect 13537 2546 13603 2549
rect 22921 2546 22987 2549
rect 11881 2544 13603 2546
rect 11881 2488 11886 2544
rect 11942 2488 13542 2544
rect 13598 2488 13603 2544
rect 11881 2486 13603 2488
rect 11881 2483 11947 2486
rect 13537 2483 13603 2486
rect 13678 2544 22987 2546
rect 13678 2488 22926 2544
rect 22982 2488 22987 2544
rect 13678 2486 22987 2488
rect 10961 2410 11027 2413
rect 2822 2408 11027 2410
rect 2822 2352 10966 2408
rect 11022 2352 11027 2408
rect 2822 2350 11027 2352
rect 0 2274 120 2304
rect 2822 2274 2882 2350
rect 10961 2347 11027 2350
rect 11237 2410 11303 2413
rect 13678 2410 13738 2486
rect 22921 2483 22987 2486
rect 24117 2546 24183 2549
rect 32857 2546 32923 2549
rect 24117 2544 32923 2546
rect 24117 2488 24122 2544
rect 24178 2488 32862 2544
rect 32918 2488 32923 2544
rect 24117 2486 32923 2488
rect 24117 2483 24183 2486
rect 32857 2483 32923 2486
rect 38377 2546 38443 2549
rect 39808 2546 39928 2576
rect 38377 2544 39928 2546
rect 38377 2488 38382 2544
rect 38438 2488 39928 2544
rect 38377 2486 39928 2488
rect 38377 2483 38443 2486
rect 39808 2456 39928 2486
rect 11237 2408 13738 2410
rect 11237 2352 11242 2408
rect 11298 2352 13738 2408
rect 11237 2350 13738 2352
rect 15469 2410 15535 2413
rect 29729 2410 29795 2413
rect 15469 2408 29795 2410
rect 15469 2352 15474 2408
rect 15530 2352 29734 2408
rect 29790 2352 29795 2408
rect 15469 2350 29795 2352
rect 11237 2347 11303 2350
rect 15469 2347 15535 2350
rect 29729 2347 29795 2350
rect 0 2214 2882 2274
rect 38009 2274 38075 2277
rect 39808 2274 39928 2304
rect 38009 2272 39928 2274
rect 38009 2216 38014 2272
rect 38070 2216 39928 2272
rect 38009 2214 39928 2216
rect 0 2184 120 2214
rect 38009 2211 38075 2214
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 9006 2208 9322 2209
rect 9006 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9322 2208
rect 9006 2143 9322 2144
rect 15006 2208 15322 2209
rect 15006 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15322 2208
rect 15006 2143 15322 2144
rect 21006 2208 21322 2209
rect 21006 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21322 2208
rect 21006 2143 21322 2144
rect 27006 2208 27322 2209
rect 27006 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27322 2208
rect 27006 2143 27322 2144
rect 33006 2208 33322 2209
rect 33006 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33322 2208
rect 39808 2184 39928 2214
rect 33006 2143 33322 2144
rect 0 2002 120 2032
rect 5717 2002 5783 2005
rect 0 2000 5783 2002
rect 0 1944 5722 2000
rect 5778 1944 5783 2000
rect 0 1942 5783 1944
rect 0 1912 120 1942
rect 5717 1939 5783 1942
rect 9949 2002 10015 2005
rect 15561 2002 15627 2005
rect 9949 2000 15627 2002
rect 9949 1944 9954 2000
rect 10010 1944 15566 2000
rect 15622 1944 15627 2000
rect 9949 1942 15627 1944
rect 9949 1939 10015 1942
rect 15561 1939 15627 1942
rect 36629 2002 36695 2005
rect 39808 2002 39928 2032
rect 36629 2000 39928 2002
rect 36629 1944 36634 2000
rect 36690 1944 39928 2000
rect 36629 1942 39928 1944
rect 36629 1939 36695 1942
rect 39808 1912 39928 1942
rect 16297 1866 16363 1869
rect 28257 1866 28323 1869
rect 16297 1864 28323 1866
rect 16297 1808 16302 1864
rect 16358 1808 28262 1864
rect 28318 1808 28323 1864
rect 16297 1806 28323 1808
rect 16297 1803 16363 1806
rect 28257 1803 28323 1806
rect 0 1730 120 1760
rect 9581 1730 9647 1733
rect 0 1728 9647 1730
rect 0 1672 9586 1728
rect 9642 1672 9647 1728
rect 0 1670 9647 1672
rect 0 1640 120 1670
rect 9581 1667 9647 1670
rect 16849 1730 16915 1733
rect 24945 1730 25011 1733
rect 16849 1728 25011 1730
rect 16849 1672 16854 1728
rect 16910 1672 24950 1728
rect 25006 1672 25011 1728
rect 16849 1670 25011 1672
rect 16849 1667 16915 1670
rect 24945 1667 25011 1670
rect 37825 1730 37891 1733
rect 39808 1730 39928 1760
rect 37825 1728 39928 1730
rect 37825 1672 37830 1728
rect 37886 1672 39928 1728
rect 37825 1670 39928 1672
rect 37825 1667 37891 1670
rect 39808 1640 39928 1670
rect 11145 1594 11211 1597
rect 20529 1594 20595 1597
rect 11145 1592 20595 1594
rect 11145 1536 11150 1592
rect 11206 1536 20534 1592
rect 20590 1536 20595 1592
rect 11145 1534 20595 1536
rect 11145 1531 11211 1534
rect 20529 1531 20595 1534
rect 0 1458 120 1488
rect 5625 1458 5691 1461
rect 0 1456 5691 1458
rect 0 1400 5630 1456
rect 5686 1400 5691 1456
rect 0 1398 5691 1400
rect 0 1368 120 1398
rect 5625 1395 5691 1398
rect 22553 1458 22619 1461
rect 31477 1458 31543 1461
rect 22553 1456 31543 1458
rect 22553 1400 22558 1456
rect 22614 1400 31482 1456
rect 31538 1400 31543 1456
rect 22553 1398 31543 1400
rect 22553 1395 22619 1398
rect 31477 1395 31543 1398
rect 37181 1458 37247 1461
rect 39808 1458 39928 1488
rect 37181 1456 39928 1458
rect 37181 1400 37186 1456
rect 37242 1400 39928 1456
rect 37181 1398 39928 1400
rect 37181 1395 37247 1398
rect 39808 1368 39928 1398
rect 0 1186 120 1216
rect 20621 1186 20687 1189
rect 0 1184 20687 1186
rect 0 1128 20626 1184
rect 20682 1128 20687 1184
rect 0 1126 20687 1128
rect 0 1096 120 1126
rect 20621 1123 20687 1126
rect 37641 1186 37707 1189
rect 39808 1186 39928 1216
rect 37641 1184 39928 1186
rect 37641 1128 37646 1184
rect 37702 1128 39928 1184
rect 37641 1126 39928 1128
rect 37641 1123 37707 1126
rect 39808 1096 39928 1126
rect 13261 642 13327 645
rect 24209 642 24275 645
rect 13261 640 24275 642
rect 13261 584 13266 640
rect 13322 584 24214 640
rect 24270 584 24275 640
rect 13261 582 24275 584
rect 13261 579 13327 582
rect 24209 579 24275 582
rect 13537 506 13603 509
rect 26141 506 26207 509
rect 13537 504 26207 506
rect 13537 448 13542 504
rect 13598 448 26146 504
rect 26202 448 26207 504
rect 13537 446 26207 448
rect 13537 443 13603 446
rect 26141 443 26207 446
rect 12709 370 12775 373
rect 25037 370 25103 373
rect 12709 368 25103 370
rect 12709 312 12714 368
rect 12770 312 25042 368
rect 25098 312 25103 368
rect 12709 310 25103 312
rect 12709 307 12775 310
rect 25037 307 25103 310
rect 14917 234 14983 237
rect 29361 234 29427 237
rect 14917 232 29427 234
rect 14917 176 14922 232
rect 14978 176 29366 232
rect 29422 176 29427 232
rect 14917 174 29427 176
rect 14917 171 14983 174
rect 29361 171 29427 174
rect 14641 98 14707 101
rect 30833 98 30899 101
rect 14641 96 30899 98
rect 14641 40 14646 96
rect 14702 40 30838 96
rect 30894 40 30899 96
rect 14641 38 30899 40
rect 14641 35 14707 38
rect 30833 35 30899 38
<< via3 >>
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 9172 8732 9236 8736
rect 9172 8676 9176 8732
rect 9176 8676 9232 8732
rect 9232 8676 9236 8732
rect 9172 8672 9236 8676
rect 9252 8732 9316 8736
rect 9252 8676 9256 8732
rect 9256 8676 9312 8732
rect 9312 8676 9316 8732
rect 9252 8672 9316 8676
rect 15012 8732 15076 8736
rect 15012 8676 15016 8732
rect 15016 8676 15072 8732
rect 15072 8676 15076 8732
rect 15012 8672 15076 8676
rect 15092 8732 15156 8736
rect 15092 8676 15096 8732
rect 15096 8676 15152 8732
rect 15152 8676 15156 8732
rect 15092 8672 15156 8676
rect 15172 8732 15236 8736
rect 15172 8676 15176 8732
rect 15176 8676 15232 8732
rect 15232 8676 15236 8732
rect 15172 8672 15236 8676
rect 15252 8732 15316 8736
rect 15252 8676 15256 8732
rect 15256 8676 15312 8732
rect 15312 8676 15316 8732
rect 15252 8672 15316 8676
rect 21012 8732 21076 8736
rect 21012 8676 21016 8732
rect 21016 8676 21072 8732
rect 21072 8676 21076 8732
rect 21012 8672 21076 8676
rect 21092 8732 21156 8736
rect 21092 8676 21096 8732
rect 21096 8676 21152 8732
rect 21152 8676 21156 8732
rect 21092 8672 21156 8676
rect 21172 8732 21236 8736
rect 21172 8676 21176 8732
rect 21176 8676 21232 8732
rect 21232 8676 21236 8732
rect 21172 8672 21236 8676
rect 21252 8732 21316 8736
rect 21252 8676 21256 8732
rect 21256 8676 21312 8732
rect 21312 8676 21316 8732
rect 21252 8672 21316 8676
rect 27012 8732 27076 8736
rect 27012 8676 27016 8732
rect 27016 8676 27072 8732
rect 27072 8676 27076 8732
rect 27012 8672 27076 8676
rect 27092 8732 27156 8736
rect 27092 8676 27096 8732
rect 27096 8676 27152 8732
rect 27152 8676 27156 8732
rect 27092 8672 27156 8676
rect 27172 8732 27236 8736
rect 27172 8676 27176 8732
rect 27176 8676 27232 8732
rect 27232 8676 27236 8732
rect 27172 8672 27236 8676
rect 27252 8732 27316 8736
rect 27252 8676 27256 8732
rect 27256 8676 27312 8732
rect 27312 8676 27316 8732
rect 27252 8672 27316 8676
rect 33012 8732 33076 8736
rect 33012 8676 33016 8732
rect 33016 8676 33072 8732
rect 33072 8676 33076 8732
rect 33012 8672 33076 8676
rect 33092 8732 33156 8736
rect 33092 8676 33096 8732
rect 33096 8676 33152 8732
rect 33152 8676 33156 8732
rect 33092 8672 33156 8676
rect 33172 8732 33236 8736
rect 33172 8676 33176 8732
rect 33176 8676 33232 8732
rect 33232 8676 33236 8732
rect 33172 8672 33236 8676
rect 33252 8732 33316 8736
rect 33252 8676 33256 8732
rect 33256 8676 33312 8732
rect 33312 8676 33316 8732
rect 33252 8672 33316 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 13952 8188 14016 8192
rect 13952 8132 13956 8188
rect 13956 8132 14012 8188
rect 14012 8132 14016 8188
rect 13952 8128 14016 8132
rect 14032 8188 14096 8192
rect 14032 8132 14036 8188
rect 14036 8132 14092 8188
rect 14092 8132 14096 8188
rect 14032 8128 14096 8132
rect 14112 8188 14176 8192
rect 14112 8132 14116 8188
rect 14116 8132 14172 8188
rect 14172 8132 14176 8188
rect 14112 8128 14176 8132
rect 14192 8188 14256 8192
rect 14192 8132 14196 8188
rect 14196 8132 14252 8188
rect 14252 8132 14256 8188
rect 14192 8128 14256 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 20192 8188 20256 8192
rect 20192 8132 20196 8188
rect 20196 8132 20252 8188
rect 20252 8132 20256 8188
rect 20192 8128 20256 8132
rect 25952 8188 26016 8192
rect 25952 8132 25956 8188
rect 25956 8132 26012 8188
rect 26012 8132 26016 8188
rect 25952 8128 26016 8132
rect 26032 8188 26096 8192
rect 26032 8132 26036 8188
rect 26036 8132 26092 8188
rect 26092 8132 26096 8188
rect 26032 8128 26096 8132
rect 26112 8188 26176 8192
rect 26112 8132 26116 8188
rect 26116 8132 26172 8188
rect 26172 8132 26176 8188
rect 26112 8128 26176 8132
rect 26192 8188 26256 8192
rect 26192 8132 26196 8188
rect 26196 8132 26252 8188
rect 26252 8132 26256 8188
rect 26192 8128 26256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 37952 8188 38016 8192
rect 37952 8132 37956 8188
rect 37956 8132 38012 8188
rect 38012 8132 38016 8188
rect 37952 8128 38016 8132
rect 38032 8188 38096 8192
rect 38032 8132 38036 8188
rect 38036 8132 38092 8188
rect 38092 8132 38096 8188
rect 38032 8128 38096 8132
rect 38112 8188 38176 8192
rect 38112 8132 38116 8188
rect 38116 8132 38172 8188
rect 38172 8132 38176 8188
rect 38112 8128 38176 8132
rect 38192 8188 38256 8192
rect 38192 8132 38196 8188
rect 38196 8132 38252 8188
rect 38252 8132 38256 8188
rect 38192 8128 38256 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 9172 7644 9236 7648
rect 9172 7588 9176 7644
rect 9176 7588 9232 7644
rect 9232 7588 9236 7644
rect 9172 7584 9236 7588
rect 9252 7644 9316 7648
rect 9252 7588 9256 7644
rect 9256 7588 9312 7644
rect 9312 7588 9316 7644
rect 9252 7584 9316 7588
rect 15012 7644 15076 7648
rect 15012 7588 15016 7644
rect 15016 7588 15072 7644
rect 15072 7588 15076 7644
rect 15012 7584 15076 7588
rect 15092 7644 15156 7648
rect 15092 7588 15096 7644
rect 15096 7588 15152 7644
rect 15152 7588 15156 7644
rect 15092 7584 15156 7588
rect 15172 7644 15236 7648
rect 15172 7588 15176 7644
rect 15176 7588 15232 7644
rect 15232 7588 15236 7644
rect 15172 7584 15236 7588
rect 15252 7644 15316 7648
rect 15252 7588 15256 7644
rect 15256 7588 15312 7644
rect 15312 7588 15316 7644
rect 15252 7584 15316 7588
rect 21012 7644 21076 7648
rect 21012 7588 21016 7644
rect 21016 7588 21072 7644
rect 21072 7588 21076 7644
rect 21012 7584 21076 7588
rect 21092 7644 21156 7648
rect 21092 7588 21096 7644
rect 21096 7588 21152 7644
rect 21152 7588 21156 7644
rect 21092 7584 21156 7588
rect 21172 7644 21236 7648
rect 21172 7588 21176 7644
rect 21176 7588 21232 7644
rect 21232 7588 21236 7644
rect 21172 7584 21236 7588
rect 21252 7644 21316 7648
rect 21252 7588 21256 7644
rect 21256 7588 21312 7644
rect 21312 7588 21316 7644
rect 21252 7584 21316 7588
rect 27012 7644 27076 7648
rect 27012 7588 27016 7644
rect 27016 7588 27072 7644
rect 27072 7588 27076 7644
rect 27012 7584 27076 7588
rect 27092 7644 27156 7648
rect 27092 7588 27096 7644
rect 27096 7588 27152 7644
rect 27152 7588 27156 7644
rect 27092 7584 27156 7588
rect 27172 7644 27236 7648
rect 27172 7588 27176 7644
rect 27176 7588 27232 7644
rect 27232 7588 27236 7644
rect 27172 7584 27236 7588
rect 27252 7644 27316 7648
rect 27252 7588 27256 7644
rect 27256 7588 27312 7644
rect 27312 7588 27316 7644
rect 27252 7584 27316 7588
rect 33012 7644 33076 7648
rect 33012 7588 33016 7644
rect 33016 7588 33072 7644
rect 33072 7588 33076 7644
rect 33012 7584 33076 7588
rect 33092 7644 33156 7648
rect 33092 7588 33096 7644
rect 33096 7588 33152 7644
rect 33152 7588 33156 7644
rect 33092 7584 33156 7588
rect 33172 7644 33236 7648
rect 33172 7588 33176 7644
rect 33176 7588 33232 7644
rect 33232 7588 33236 7644
rect 33172 7584 33236 7588
rect 33252 7644 33316 7648
rect 33252 7588 33256 7644
rect 33256 7588 33312 7644
rect 33312 7588 33316 7644
rect 33252 7584 33316 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 13952 7100 14016 7104
rect 13952 7044 13956 7100
rect 13956 7044 14012 7100
rect 14012 7044 14016 7100
rect 13952 7040 14016 7044
rect 14032 7100 14096 7104
rect 14032 7044 14036 7100
rect 14036 7044 14092 7100
rect 14092 7044 14096 7100
rect 14032 7040 14096 7044
rect 14112 7100 14176 7104
rect 14112 7044 14116 7100
rect 14116 7044 14172 7100
rect 14172 7044 14176 7100
rect 14112 7040 14176 7044
rect 14192 7100 14256 7104
rect 14192 7044 14196 7100
rect 14196 7044 14252 7100
rect 14252 7044 14256 7100
rect 14192 7040 14256 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 20192 7100 20256 7104
rect 20192 7044 20196 7100
rect 20196 7044 20252 7100
rect 20252 7044 20256 7100
rect 20192 7040 20256 7044
rect 25952 7100 26016 7104
rect 25952 7044 25956 7100
rect 25956 7044 26012 7100
rect 26012 7044 26016 7100
rect 25952 7040 26016 7044
rect 26032 7100 26096 7104
rect 26032 7044 26036 7100
rect 26036 7044 26092 7100
rect 26092 7044 26096 7100
rect 26032 7040 26096 7044
rect 26112 7100 26176 7104
rect 26112 7044 26116 7100
rect 26116 7044 26172 7100
rect 26172 7044 26176 7100
rect 26112 7040 26176 7044
rect 26192 7100 26256 7104
rect 26192 7044 26196 7100
rect 26196 7044 26252 7100
rect 26252 7044 26256 7100
rect 26192 7040 26256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 37952 7100 38016 7104
rect 37952 7044 37956 7100
rect 37956 7044 38012 7100
rect 38012 7044 38016 7100
rect 37952 7040 38016 7044
rect 38032 7100 38096 7104
rect 38032 7044 38036 7100
rect 38036 7044 38092 7100
rect 38092 7044 38096 7100
rect 38032 7040 38096 7044
rect 38112 7100 38176 7104
rect 38112 7044 38116 7100
rect 38116 7044 38172 7100
rect 38172 7044 38176 7100
rect 38112 7040 38176 7044
rect 38192 7100 38256 7104
rect 38192 7044 38196 7100
rect 38196 7044 38252 7100
rect 38252 7044 38256 7100
rect 38192 7040 38256 7044
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 9172 6556 9236 6560
rect 9172 6500 9176 6556
rect 9176 6500 9232 6556
rect 9232 6500 9236 6556
rect 9172 6496 9236 6500
rect 9252 6556 9316 6560
rect 9252 6500 9256 6556
rect 9256 6500 9312 6556
rect 9312 6500 9316 6556
rect 9252 6496 9316 6500
rect 15012 6556 15076 6560
rect 15012 6500 15016 6556
rect 15016 6500 15072 6556
rect 15072 6500 15076 6556
rect 15012 6496 15076 6500
rect 15092 6556 15156 6560
rect 15092 6500 15096 6556
rect 15096 6500 15152 6556
rect 15152 6500 15156 6556
rect 15092 6496 15156 6500
rect 15172 6556 15236 6560
rect 15172 6500 15176 6556
rect 15176 6500 15232 6556
rect 15232 6500 15236 6556
rect 15172 6496 15236 6500
rect 15252 6556 15316 6560
rect 15252 6500 15256 6556
rect 15256 6500 15312 6556
rect 15312 6500 15316 6556
rect 15252 6496 15316 6500
rect 21012 6556 21076 6560
rect 21012 6500 21016 6556
rect 21016 6500 21072 6556
rect 21072 6500 21076 6556
rect 21012 6496 21076 6500
rect 21092 6556 21156 6560
rect 21092 6500 21096 6556
rect 21096 6500 21152 6556
rect 21152 6500 21156 6556
rect 21092 6496 21156 6500
rect 21172 6556 21236 6560
rect 21172 6500 21176 6556
rect 21176 6500 21232 6556
rect 21232 6500 21236 6556
rect 21172 6496 21236 6500
rect 21252 6556 21316 6560
rect 21252 6500 21256 6556
rect 21256 6500 21312 6556
rect 21312 6500 21316 6556
rect 21252 6496 21316 6500
rect 27012 6556 27076 6560
rect 27012 6500 27016 6556
rect 27016 6500 27072 6556
rect 27072 6500 27076 6556
rect 27012 6496 27076 6500
rect 27092 6556 27156 6560
rect 27092 6500 27096 6556
rect 27096 6500 27152 6556
rect 27152 6500 27156 6556
rect 27092 6496 27156 6500
rect 27172 6556 27236 6560
rect 27172 6500 27176 6556
rect 27176 6500 27232 6556
rect 27232 6500 27236 6556
rect 27172 6496 27236 6500
rect 27252 6556 27316 6560
rect 27252 6500 27256 6556
rect 27256 6500 27312 6556
rect 27312 6500 27316 6556
rect 27252 6496 27316 6500
rect 33012 6556 33076 6560
rect 33012 6500 33016 6556
rect 33016 6500 33072 6556
rect 33072 6500 33076 6556
rect 33012 6496 33076 6500
rect 33092 6556 33156 6560
rect 33092 6500 33096 6556
rect 33096 6500 33152 6556
rect 33152 6500 33156 6556
rect 33092 6496 33156 6500
rect 33172 6556 33236 6560
rect 33172 6500 33176 6556
rect 33176 6500 33232 6556
rect 33232 6500 33236 6556
rect 33172 6496 33236 6500
rect 33252 6556 33316 6560
rect 33252 6500 33256 6556
rect 33256 6500 33312 6556
rect 33312 6500 33316 6556
rect 33252 6496 33316 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 13952 6012 14016 6016
rect 13952 5956 13956 6012
rect 13956 5956 14012 6012
rect 14012 5956 14016 6012
rect 13952 5952 14016 5956
rect 14032 6012 14096 6016
rect 14032 5956 14036 6012
rect 14036 5956 14092 6012
rect 14092 5956 14096 6012
rect 14032 5952 14096 5956
rect 14112 6012 14176 6016
rect 14112 5956 14116 6012
rect 14116 5956 14172 6012
rect 14172 5956 14176 6012
rect 14112 5952 14176 5956
rect 14192 6012 14256 6016
rect 14192 5956 14196 6012
rect 14196 5956 14252 6012
rect 14252 5956 14256 6012
rect 14192 5952 14256 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 20192 6012 20256 6016
rect 20192 5956 20196 6012
rect 20196 5956 20252 6012
rect 20252 5956 20256 6012
rect 20192 5952 20256 5956
rect 25952 6012 26016 6016
rect 25952 5956 25956 6012
rect 25956 5956 26012 6012
rect 26012 5956 26016 6012
rect 25952 5952 26016 5956
rect 26032 6012 26096 6016
rect 26032 5956 26036 6012
rect 26036 5956 26092 6012
rect 26092 5956 26096 6012
rect 26032 5952 26096 5956
rect 26112 6012 26176 6016
rect 26112 5956 26116 6012
rect 26116 5956 26172 6012
rect 26172 5956 26176 6012
rect 26112 5952 26176 5956
rect 26192 6012 26256 6016
rect 26192 5956 26196 6012
rect 26196 5956 26252 6012
rect 26252 5956 26256 6012
rect 26192 5952 26256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 37952 6012 38016 6016
rect 37952 5956 37956 6012
rect 37956 5956 38012 6012
rect 38012 5956 38016 6012
rect 37952 5952 38016 5956
rect 38032 6012 38096 6016
rect 38032 5956 38036 6012
rect 38036 5956 38092 6012
rect 38092 5956 38096 6012
rect 38032 5952 38096 5956
rect 38112 6012 38176 6016
rect 38112 5956 38116 6012
rect 38116 5956 38172 6012
rect 38172 5956 38176 6012
rect 38112 5952 38176 5956
rect 38192 6012 38256 6016
rect 38192 5956 38196 6012
rect 38196 5956 38252 6012
rect 38252 5956 38256 6012
rect 38192 5952 38256 5956
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 9172 5468 9236 5472
rect 9172 5412 9176 5468
rect 9176 5412 9232 5468
rect 9232 5412 9236 5468
rect 9172 5408 9236 5412
rect 9252 5468 9316 5472
rect 9252 5412 9256 5468
rect 9256 5412 9312 5468
rect 9312 5412 9316 5468
rect 9252 5408 9316 5412
rect 15012 5468 15076 5472
rect 15012 5412 15016 5468
rect 15016 5412 15072 5468
rect 15072 5412 15076 5468
rect 15012 5408 15076 5412
rect 15092 5468 15156 5472
rect 15092 5412 15096 5468
rect 15096 5412 15152 5468
rect 15152 5412 15156 5468
rect 15092 5408 15156 5412
rect 15172 5468 15236 5472
rect 15172 5412 15176 5468
rect 15176 5412 15232 5468
rect 15232 5412 15236 5468
rect 15172 5408 15236 5412
rect 15252 5468 15316 5472
rect 15252 5412 15256 5468
rect 15256 5412 15312 5468
rect 15312 5412 15316 5468
rect 15252 5408 15316 5412
rect 21012 5468 21076 5472
rect 21012 5412 21016 5468
rect 21016 5412 21072 5468
rect 21072 5412 21076 5468
rect 21012 5408 21076 5412
rect 21092 5468 21156 5472
rect 21092 5412 21096 5468
rect 21096 5412 21152 5468
rect 21152 5412 21156 5468
rect 21092 5408 21156 5412
rect 21172 5468 21236 5472
rect 21172 5412 21176 5468
rect 21176 5412 21232 5468
rect 21232 5412 21236 5468
rect 21172 5408 21236 5412
rect 21252 5468 21316 5472
rect 21252 5412 21256 5468
rect 21256 5412 21312 5468
rect 21312 5412 21316 5468
rect 21252 5408 21316 5412
rect 27012 5468 27076 5472
rect 27012 5412 27016 5468
rect 27016 5412 27072 5468
rect 27072 5412 27076 5468
rect 27012 5408 27076 5412
rect 27092 5468 27156 5472
rect 27092 5412 27096 5468
rect 27096 5412 27152 5468
rect 27152 5412 27156 5468
rect 27092 5408 27156 5412
rect 27172 5468 27236 5472
rect 27172 5412 27176 5468
rect 27176 5412 27232 5468
rect 27232 5412 27236 5468
rect 27172 5408 27236 5412
rect 27252 5468 27316 5472
rect 27252 5412 27256 5468
rect 27256 5412 27312 5468
rect 27312 5412 27316 5468
rect 27252 5408 27316 5412
rect 33012 5468 33076 5472
rect 33012 5412 33016 5468
rect 33016 5412 33072 5468
rect 33072 5412 33076 5468
rect 33012 5408 33076 5412
rect 33092 5468 33156 5472
rect 33092 5412 33096 5468
rect 33096 5412 33152 5468
rect 33152 5412 33156 5468
rect 33092 5408 33156 5412
rect 33172 5468 33236 5472
rect 33172 5412 33176 5468
rect 33176 5412 33232 5468
rect 33232 5412 33236 5468
rect 33172 5408 33236 5412
rect 33252 5468 33316 5472
rect 33252 5412 33256 5468
rect 33256 5412 33312 5468
rect 33312 5412 33316 5468
rect 33252 5408 33316 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 13952 4924 14016 4928
rect 13952 4868 13956 4924
rect 13956 4868 14012 4924
rect 14012 4868 14016 4924
rect 13952 4864 14016 4868
rect 14032 4924 14096 4928
rect 14032 4868 14036 4924
rect 14036 4868 14092 4924
rect 14092 4868 14096 4924
rect 14032 4864 14096 4868
rect 14112 4924 14176 4928
rect 14112 4868 14116 4924
rect 14116 4868 14172 4924
rect 14172 4868 14176 4924
rect 14112 4864 14176 4868
rect 14192 4924 14256 4928
rect 14192 4868 14196 4924
rect 14196 4868 14252 4924
rect 14252 4868 14256 4924
rect 14192 4864 14256 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 20192 4924 20256 4928
rect 20192 4868 20196 4924
rect 20196 4868 20252 4924
rect 20252 4868 20256 4924
rect 20192 4864 20256 4868
rect 25952 4924 26016 4928
rect 25952 4868 25956 4924
rect 25956 4868 26012 4924
rect 26012 4868 26016 4924
rect 25952 4864 26016 4868
rect 26032 4924 26096 4928
rect 26032 4868 26036 4924
rect 26036 4868 26092 4924
rect 26092 4868 26096 4924
rect 26032 4864 26096 4868
rect 26112 4924 26176 4928
rect 26112 4868 26116 4924
rect 26116 4868 26172 4924
rect 26172 4868 26176 4924
rect 26112 4864 26176 4868
rect 26192 4924 26256 4928
rect 26192 4868 26196 4924
rect 26196 4868 26252 4924
rect 26252 4868 26256 4924
rect 26192 4864 26256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 37952 4924 38016 4928
rect 37952 4868 37956 4924
rect 37956 4868 38012 4924
rect 38012 4868 38016 4924
rect 37952 4864 38016 4868
rect 38032 4924 38096 4928
rect 38032 4868 38036 4924
rect 38036 4868 38092 4924
rect 38092 4868 38096 4924
rect 38032 4864 38096 4868
rect 38112 4924 38176 4928
rect 38112 4868 38116 4924
rect 38116 4868 38172 4924
rect 38172 4868 38176 4924
rect 38112 4864 38176 4868
rect 38192 4924 38256 4928
rect 38192 4868 38196 4924
rect 38196 4868 38252 4924
rect 38252 4868 38256 4924
rect 38192 4864 38256 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 9172 4380 9236 4384
rect 9172 4324 9176 4380
rect 9176 4324 9232 4380
rect 9232 4324 9236 4380
rect 9172 4320 9236 4324
rect 9252 4380 9316 4384
rect 9252 4324 9256 4380
rect 9256 4324 9312 4380
rect 9312 4324 9316 4380
rect 9252 4320 9316 4324
rect 15012 4380 15076 4384
rect 15012 4324 15016 4380
rect 15016 4324 15072 4380
rect 15072 4324 15076 4380
rect 15012 4320 15076 4324
rect 15092 4380 15156 4384
rect 15092 4324 15096 4380
rect 15096 4324 15152 4380
rect 15152 4324 15156 4380
rect 15092 4320 15156 4324
rect 15172 4380 15236 4384
rect 15172 4324 15176 4380
rect 15176 4324 15232 4380
rect 15232 4324 15236 4380
rect 15172 4320 15236 4324
rect 15252 4380 15316 4384
rect 15252 4324 15256 4380
rect 15256 4324 15312 4380
rect 15312 4324 15316 4380
rect 15252 4320 15316 4324
rect 21012 4380 21076 4384
rect 21012 4324 21016 4380
rect 21016 4324 21072 4380
rect 21072 4324 21076 4380
rect 21012 4320 21076 4324
rect 21092 4380 21156 4384
rect 21092 4324 21096 4380
rect 21096 4324 21152 4380
rect 21152 4324 21156 4380
rect 21092 4320 21156 4324
rect 21172 4380 21236 4384
rect 21172 4324 21176 4380
rect 21176 4324 21232 4380
rect 21232 4324 21236 4380
rect 21172 4320 21236 4324
rect 21252 4380 21316 4384
rect 21252 4324 21256 4380
rect 21256 4324 21312 4380
rect 21312 4324 21316 4380
rect 21252 4320 21316 4324
rect 27012 4380 27076 4384
rect 27012 4324 27016 4380
rect 27016 4324 27072 4380
rect 27072 4324 27076 4380
rect 27012 4320 27076 4324
rect 27092 4380 27156 4384
rect 27092 4324 27096 4380
rect 27096 4324 27152 4380
rect 27152 4324 27156 4380
rect 27092 4320 27156 4324
rect 27172 4380 27236 4384
rect 27172 4324 27176 4380
rect 27176 4324 27232 4380
rect 27232 4324 27236 4380
rect 27172 4320 27236 4324
rect 27252 4380 27316 4384
rect 27252 4324 27256 4380
rect 27256 4324 27312 4380
rect 27312 4324 27316 4380
rect 27252 4320 27316 4324
rect 33012 4380 33076 4384
rect 33012 4324 33016 4380
rect 33016 4324 33072 4380
rect 33072 4324 33076 4380
rect 33012 4320 33076 4324
rect 33092 4380 33156 4384
rect 33092 4324 33096 4380
rect 33096 4324 33152 4380
rect 33152 4324 33156 4380
rect 33092 4320 33156 4324
rect 33172 4380 33236 4384
rect 33172 4324 33176 4380
rect 33176 4324 33232 4380
rect 33232 4324 33236 4380
rect 33172 4320 33236 4324
rect 33252 4380 33316 4384
rect 33252 4324 33256 4380
rect 33256 4324 33312 4380
rect 33312 4324 33316 4380
rect 33252 4320 33316 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 13952 3836 14016 3840
rect 13952 3780 13956 3836
rect 13956 3780 14012 3836
rect 14012 3780 14016 3836
rect 13952 3776 14016 3780
rect 14032 3836 14096 3840
rect 14032 3780 14036 3836
rect 14036 3780 14092 3836
rect 14092 3780 14096 3836
rect 14032 3776 14096 3780
rect 14112 3836 14176 3840
rect 14112 3780 14116 3836
rect 14116 3780 14172 3836
rect 14172 3780 14176 3836
rect 14112 3776 14176 3780
rect 14192 3836 14256 3840
rect 14192 3780 14196 3836
rect 14196 3780 14252 3836
rect 14252 3780 14256 3836
rect 14192 3776 14256 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 20192 3836 20256 3840
rect 20192 3780 20196 3836
rect 20196 3780 20252 3836
rect 20252 3780 20256 3836
rect 20192 3776 20256 3780
rect 25952 3836 26016 3840
rect 25952 3780 25956 3836
rect 25956 3780 26012 3836
rect 26012 3780 26016 3836
rect 25952 3776 26016 3780
rect 26032 3836 26096 3840
rect 26032 3780 26036 3836
rect 26036 3780 26092 3836
rect 26092 3780 26096 3836
rect 26032 3776 26096 3780
rect 26112 3836 26176 3840
rect 26112 3780 26116 3836
rect 26116 3780 26172 3836
rect 26172 3780 26176 3836
rect 26112 3776 26176 3780
rect 26192 3836 26256 3840
rect 26192 3780 26196 3836
rect 26196 3780 26252 3836
rect 26252 3780 26256 3836
rect 26192 3776 26256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 37952 3836 38016 3840
rect 37952 3780 37956 3836
rect 37956 3780 38012 3836
rect 38012 3780 38016 3836
rect 37952 3776 38016 3780
rect 38032 3836 38096 3840
rect 38032 3780 38036 3836
rect 38036 3780 38092 3836
rect 38092 3780 38096 3836
rect 38032 3776 38096 3780
rect 38112 3836 38176 3840
rect 38112 3780 38116 3836
rect 38116 3780 38172 3836
rect 38172 3780 38176 3836
rect 38112 3776 38176 3780
rect 38192 3836 38256 3840
rect 38192 3780 38196 3836
rect 38196 3780 38252 3836
rect 38252 3780 38256 3836
rect 38192 3776 38256 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 9172 3292 9236 3296
rect 9172 3236 9176 3292
rect 9176 3236 9232 3292
rect 9232 3236 9236 3292
rect 9172 3232 9236 3236
rect 9252 3292 9316 3296
rect 9252 3236 9256 3292
rect 9256 3236 9312 3292
rect 9312 3236 9316 3292
rect 9252 3232 9316 3236
rect 15012 3292 15076 3296
rect 15012 3236 15016 3292
rect 15016 3236 15072 3292
rect 15072 3236 15076 3292
rect 15012 3232 15076 3236
rect 15092 3292 15156 3296
rect 15092 3236 15096 3292
rect 15096 3236 15152 3292
rect 15152 3236 15156 3292
rect 15092 3232 15156 3236
rect 15172 3292 15236 3296
rect 15172 3236 15176 3292
rect 15176 3236 15232 3292
rect 15232 3236 15236 3292
rect 15172 3232 15236 3236
rect 15252 3292 15316 3296
rect 15252 3236 15256 3292
rect 15256 3236 15312 3292
rect 15312 3236 15316 3292
rect 15252 3232 15316 3236
rect 21012 3292 21076 3296
rect 21012 3236 21016 3292
rect 21016 3236 21072 3292
rect 21072 3236 21076 3292
rect 21012 3232 21076 3236
rect 21092 3292 21156 3296
rect 21092 3236 21096 3292
rect 21096 3236 21152 3292
rect 21152 3236 21156 3292
rect 21092 3232 21156 3236
rect 21172 3292 21236 3296
rect 21172 3236 21176 3292
rect 21176 3236 21232 3292
rect 21232 3236 21236 3292
rect 21172 3232 21236 3236
rect 21252 3292 21316 3296
rect 21252 3236 21256 3292
rect 21256 3236 21312 3292
rect 21312 3236 21316 3292
rect 21252 3232 21316 3236
rect 27012 3292 27076 3296
rect 27012 3236 27016 3292
rect 27016 3236 27072 3292
rect 27072 3236 27076 3292
rect 27012 3232 27076 3236
rect 27092 3292 27156 3296
rect 27092 3236 27096 3292
rect 27096 3236 27152 3292
rect 27152 3236 27156 3292
rect 27092 3232 27156 3236
rect 27172 3292 27236 3296
rect 27172 3236 27176 3292
rect 27176 3236 27232 3292
rect 27232 3236 27236 3292
rect 27172 3232 27236 3236
rect 27252 3292 27316 3296
rect 27252 3236 27256 3292
rect 27256 3236 27312 3292
rect 27312 3236 27316 3292
rect 27252 3232 27316 3236
rect 33012 3292 33076 3296
rect 33012 3236 33016 3292
rect 33016 3236 33072 3292
rect 33072 3236 33076 3292
rect 33012 3232 33076 3236
rect 33092 3292 33156 3296
rect 33092 3236 33096 3292
rect 33096 3236 33152 3292
rect 33152 3236 33156 3292
rect 33092 3232 33156 3236
rect 33172 3292 33236 3296
rect 33172 3236 33176 3292
rect 33176 3236 33232 3292
rect 33232 3236 33236 3292
rect 33172 3232 33236 3236
rect 33252 3292 33316 3296
rect 33252 3236 33256 3292
rect 33256 3236 33312 3292
rect 33312 3236 33316 3292
rect 33252 3232 33316 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 13952 2748 14016 2752
rect 13952 2692 13956 2748
rect 13956 2692 14012 2748
rect 14012 2692 14016 2748
rect 13952 2688 14016 2692
rect 14032 2748 14096 2752
rect 14032 2692 14036 2748
rect 14036 2692 14092 2748
rect 14092 2692 14096 2748
rect 14032 2688 14096 2692
rect 14112 2748 14176 2752
rect 14112 2692 14116 2748
rect 14116 2692 14172 2748
rect 14172 2692 14176 2748
rect 14112 2688 14176 2692
rect 14192 2748 14256 2752
rect 14192 2692 14196 2748
rect 14196 2692 14252 2748
rect 14252 2692 14256 2748
rect 14192 2688 14256 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 20192 2748 20256 2752
rect 20192 2692 20196 2748
rect 20196 2692 20252 2748
rect 20252 2692 20256 2748
rect 20192 2688 20256 2692
rect 25952 2748 26016 2752
rect 25952 2692 25956 2748
rect 25956 2692 26012 2748
rect 26012 2692 26016 2748
rect 25952 2688 26016 2692
rect 26032 2748 26096 2752
rect 26032 2692 26036 2748
rect 26036 2692 26092 2748
rect 26092 2692 26096 2748
rect 26032 2688 26096 2692
rect 26112 2748 26176 2752
rect 26112 2692 26116 2748
rect 26116 2692 26172 2748
rect 26172 2692 26176 2748
rect 26112 2688 26176 2692
rect 26192 2748 26256 2752
rect 26192 2692 26196 2748
rect 26196 2692 26252 2748
rect 26252 2692 26256 2748
rect 26192 2688 26256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 37952 2748 38016 2752
rect 37952 2692 37956 2748
rect 37956 2692 38012 2748
rect 38012 2692 38016 2748
rect 37952 2688 38016 2692
rect 38032 2748 38096 2752
rect 38032 2692 38036 2748
rect 38036 2692 38092 2748
rect 38092 2692 38096 2748
rect 38032 2688 38096 2692
rect 38112 2748 38176 2752
rect 38112 2692 38116 2748
rect 38116 2692 38172 2748
rect 38172 2692 38176 2748
rect 38112 2688 38176 2692
rect 38192 2748 38256 2752
rect 38192 2692 38196 2748
rect 38196 2692 38252 2748
rect 38252 2692 38256 2748
rect 38192 2688 38256 2692
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 9172 2204 9236 2208
rect 9172 2148 9176 2204
rect 9176 2148 9232 2204
rect 9232 2148 9236 2204
rect 9172 2144 9236 2148
rect 9252 2204 9316 2208
rect 9252 2148 9256 2204
rect 9256 2148 9312 2204
rect 9312 2148 9316 2204
rect 9252 2144 9316 2148
rect 15012 2204 15076 2208
rect 15012 2148 15016 2204
rect 15016 2148 15072 2204
rect 15072 2148 15076 2204
rect 15012 2144 15076 2148
rect 15092 2204 15156 2208
rect 15092 2148 15096 2204
rect 15096 2148 15152 2204
rect 15152 2148 15156 2204
rect 15092 2144 15156 2148
rect 15172 2204 15236 2208
rect 15172 2148 15176 2204
rect 15176 2148 15232 2204
rect 15232 2148 15236 2204
rect 15172 2144 15236 2148
rect 15252 2204 15316 2208
rect 15252 2148 15256 2204
rect 15256 2148 15312 2204
rect 15312 2148 15316 2204
rect 15252 2144 15316 2148
rect 21012 2204 21076 2208
rect 21012 2148 21016 2204
rect 21016 2148 21072 2204
rect 21072 2148 21076 2204
rect 21012 2144 21076 2148
rect 21092 2204 21156 2208
rect 21092 2148 21096 2204
rect 21096 2148 21152 2204
rect 21152 2148 21156 2204
rect 21092 2144 21156 2148
rect 21172 2204 21236 2208
rect 21172 2148 21176 2204
rect 21176 2148 21232 2204
rect 21232 2148 21236 2204
rect 21172 2144 21236 2148
rect 21252 2204 21316 2208
rect 21252 2148 21256 2204
rect 21256 2148 21312 2204
rect 21312 2148 21316 2204
rect 21252 2144 21316 2148
rect 27012 2204 27076 2208
rect 27012 2148 27016 2204
rect 27016 2148 27072 2204
rect 27072 2148 27076 2204
rect 27012 2144 27076 2148
rect 27092 2204 27156 2208
rect 27092 2148 27096 2204
rect 27096 2148 27152 2204
rect 27152 2148 27156 2204
rect 27092 2144 27156 2148
rect 27172 2204 27236 2208
rect 27172 2148 27176 2204
rect 27176 2148 27232 2204
rect 27232 2148 27236 2204
rect 27172 2144 27236 2148
rect 27252 2204 27316 2208
rect 27252 2148 27256 2204
rect 27256 2148 27312 2204
rect 27312 2148 27316 2204
rect 27252 2144 27316 2148
rect 33012 2204 33076 2208
rect 33012 2148 33016 2204
rect 33016 2148 33072 2204
rect 33072 2148 33076 2204
rect 33012 2144 33076 2148
rect 33092 2204 33156 2208
rect 33092 2148 33096 2204
rect 33096 2148 33152 2204
rect 33152 2148 33156 2204
rect 33092 2144 33156 2148
rect 33172 2204 33236 2208
rect 33172 2148 33176 2204
rect 33176 2148 33232 2204
rect 33232 2148 33236 2204
rect 33172 2144 33236 2148
rect 33252 2204 33316 2208
rect 33252 2148 33256 2204
rect 33256 2148 33312 2204
rect 33312 2148 33316 2204
rect 33252 2144 33316 2148
<< metal4 >>
rect 1944 8192 2264 11152
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 0 2264 2688
rect 3004 8736 3324 11152
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 0 3324 2144
rect 7944 8192 8264 11152
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 7944 6016 8264 7040
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 4928 8264 5952
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 2752 8264 3776
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 7944 0 8264 2688
rect 9004 8736 9324 11152
rect 9004 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9324 8736
rect 9004 7648 9324 8672
rect 9004 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9324 7648
rect 9004 6560 9324 7584
rect 9004 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9324 6560
rect 9004 5472 9324 6496
rect 9004 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9324 5472
rect 9004 4384 9324 5408
rect 9004 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9324 4384
rect 9004 3296 9324 4320
rect 9004 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9324 3296
rect 9004 2208 9324 3232
rect 9004 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9324 2208
rect 9004 0 9324 2144
rect 13944 8192 14264 11152
rect 13944 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14264 8192
rect 13944 7104 14264 8128
rect 13944 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14264 7104
rect 13944 6016 14264 7040
rect 13944 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14264 6016
rect 13944 4928 14264 5952
rect 13944 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14264 4928
rect 13944 3840 14264 4864
rect 13944 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14264 3840
rect 13944 2752 14264 3776
rect 13944 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14264 2752
rect 13944 0 14264 2688
rect 15004 8736 15324 11152
rect 15004 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15324 8736
rect 15004 7648 15324 8672
rect 15004 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15324 7648
rect 15004 6560 15324 7584
rect 15004 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15324 6560
rect 15004 5472 15324 6496
rect 15004 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15324 5472
rect 15004 4384 15324 5408
rect 15004 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15324 4384
rect 15004 3296 15324 4320
rect 15004 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15324 3296
rect 15004 2208 15324 3232
rect 15004 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15324 2208
rect 15004 0 15324 2144
rect 19944 8192 20264 11152
rect 19944 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20264 8192
rect 19944 7104 20264 8128
rect 19944 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20264 7104
rect 19944 6016 20264 7040
rect 19944 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20264 6016
rect 19944 4928 20264 5952
rect 19944 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20264 4928
rect 19944 3840 20264 4864
rect 19944 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20264 3840
rect 19944 2752 20264 3776
rect 19944 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20264 2752
rect 19944 0 20264 2688
rect 21004 8736 21324 11152
rect 21004 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21324 8736
rect 21004 7648 21324 8672
rect 21004 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21324 7648
rect 21004 6560 21324 7584
rect 21004 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21324 6560
rect 21004 5472 21324 6496
rect 21004 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21324 5472
rect 21004 4384 21324 5408
rect 21004 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21324 4384
rect 21004 3296 21324 4320
rect 21004 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21324 3296
rect 21004 2208 21324 3232
rect 21004 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21324 2208
rect 21004 0 21324 2144
rect 25944 8192 26264 11152
rect 25944 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26264 8192
rect 25944 7104 26264 8128
rect 25944 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26264 7104
rect 25944 6016 26264 7040
rect 25944 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26264 6016
rect 25944 4928 26264 5952
rect 25944 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26264 4928
rect 25944 3840 26264 4864
rect 25944 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26264 3840
rect 25944 2752 26264 3776
rect 25944 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26264 2752
rect 25944 0 26264 2688
rect 27004 8736 27324 11152
rect 27004 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27324 8736
rect 27004 7648 27324 8672
rect 27004 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27324 7648
rect 27004 6560 27324 7584
rect 27004 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27324 6560
rect 27004 5472 27324 6496
rect 27004 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27324 5472
rect 27004 4384 27324 5408
rect 27004 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27324 4384
rect 27004 3296 27324 4320
rect 27004 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27324 3296
rect 27004 2208 27324 3232
rect 27004 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27324 2208
rect 27004 0 27324 2144
rect 31944 8192 32264 11152
rect 31944 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32264 8192
rect 31944 7104 32264 8128
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 2752 32264 3776
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 31944 0 32264 2688
rect 33004 8736 33324 11152
rect 33004 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33324 8736
rect 33004 7648 33324 8672
rect 33004 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33324 7648
rect 33004 6560 33324 7584
rect 33004 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33324 6560
rect 33004 5472 33324 6496
rect 33004 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33324 5472
rect 33004 4384 33324 5408
rect 33004 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33324 4384
rect 33004 3296 33324 4320
rect 33004 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33324 3296
rect 33004 2208 33324 3232
rect 33004 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33324 2208
rect 33004 0 33324 2144
rect 37944 8192 38264 11152
rect 37944 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38264 8192
rect 37944 7104 38264 8128
rect 37944 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38264 7104
rect 37944 6016 38264 7040
rect 37944 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38264 6016
rect 37944 4928 38264 5952
rect 37944 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38264 4928
rect 37944 3840 38264 4864
rect 37944 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38264 3840
rect 37944 2752 38264 3776
rect 37944 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38264 2752
rect 37944 0 38264 2688
use sky130_fd_sc_hd__buf_1  _000_
timestamp -3599
transform 1 0 21068 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _001_
timestamp -3599
transform 1 0 22080 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _002_
timestamp -3599
transform 1 0 22632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _003_
timestamp -3599
transform 1 0 22356 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _004_
timestamp -3599
transform 1 0 21620 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _005_
timestamp -3599
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _006_
timestamp -3599
transform 1 0 23920 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _007_
timestamp -3599
transform 1 0 23368 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _008_
timestamp -3599
transform 1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _009_
timestamp -3599
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _010_
timestamp -3599
transform 1 0 23552 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _011_
timestamp -3599
transform 1 0 23460 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _012_
timestamp -3599
transform 1 0 23000 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _013_
timestamp -3599
transform 1 0 21528 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _014_
timestamp -3599
transform 1 0 19228 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _015_
timestamp -3599
transform 1 0 19412 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _016_
timestamp -3599
transform 1 0 19964 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _017_
timestamp -3599
transform 1 0 21620 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _018_
timestamp -3599
transform 1 0 17572 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _019_
timestamp -3599
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _020_
timestamp -3599
transform 1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _021_
timestamp -3599
transform 1 0 15916 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _022_
timestamp -3599
transform 1 0 19964 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _023_
timestamp -3599
transform 1 0 15456 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _024_
timestamp -3599
transform 1 0 18584 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _025_
timestamp -3599
transform 1 0 18216 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _026_
timestamp -3599
transform 1 0 19504 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _027_
timestamp -3599
transform 1 0 17480 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _028_
timestamp -3599
transform 1 0 17204 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _029_
timestamp -3599
transform -1 0 16008 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _030_
timestamp -3599
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _031_
timestamp -3599
transform 1 0 19780 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _032_
timestamp -3599
transform -1 0 22080 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _033_
timestamp -3599
transform -1 0 19228 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _034_
timestamp -3599
transform -1 0 21620 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _035_
timestamp -3599
transform 1 0 17756 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _036_
timestamp -3599
transform -1 0 23920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _037_
timestamp -3599
transform -1 0 25484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _038_
timestamp -3599
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _039_
timestamp -3599
transform 1 0 26036 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _040_
timestamp -3599
transform 1 0 26312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _041_
timestamp -3599
transform 1 0 26312 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _042_
timestamp -3599
transform 1 0 28152 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _043_
timestamp -3599
transform 1 0 28796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _044_
timestamp -3599
transform 1 0 28060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp -3599
transform 1 0 29532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp -3599
transform 1 0 30728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _047_
timestamp -3599
transform 1 0 32844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp -3599
transform 1 0 34224 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp -3599
transform 1 0 35512 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _050_
timestamp -3599
transform 1 0 36708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _051_
timestamp -3599
transform -1 0 37260 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _052_
timestamp -3599
transform 1 0 2852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _053_
timestamp -3599
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _054_
timestamp -3599
transform 1 0 4232 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _055_
timestamp -3599
transform 1 0 5520 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _056_
timestamp -3599
transform 1 0 4416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _057_
timestamp -3599
transform 1 0 4140 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _058_
timestamp -3599
transform 1 0 4692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _059_
timestamp -3599
transform 1 0 5980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _060_
timestamp -3599
transform 1 0 7268 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _061_
timestamp -3599
transform 1 0 8372 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _062_
timestamp -3599
transform 1 0 9568 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _063_
timestamp -3599
transform 1 0 10396 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _064_
timestamp -3599
transform 1 0 7360 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _065_
timestamp -3599
transform 1 0 7636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _066_
timestamp -3599
transform 1 0 8096 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _067_
timestamp -3599
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _068_
timestamp -3599
transform 1 0 9292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _069_
timestamp -3599
transform 1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _070_
timestamp -3599
transform 1 0 10304 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _071_
timestamp -3599
transform 1 0 10948 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp -3599
transform -1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp -3599
transform -1 0 14260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _074_
timestamp -3599
transform 1 0 13524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _075_
timestamp -3599
transform 1 0 13156 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _076_
timestamp -3599
transform 1 0 12604 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _077_
timestamp -3599
transform 1 0 12880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _078_
timestamp -3599
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _079_
timestamp -3599
transform 1 0 13708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _080_
timestamp -3599
transform 1 0 14260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _081_
timestamp -3599
transform 1 0 15272 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _082_
timestamp -3599
transform 1 0 14996 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp -3599
transform -1 0 16192 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp -3599
transform -1 0 16652 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp -3599
transform -1 0 17112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp -3599
transform -1 0 18032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp -3599
transform -1 0 17756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp -3599
transform -1 0 27324 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp -3599
transform -1 0 27968 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp -3599
transform 1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp -3599
transform 1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp -3599
transform 1 0 29532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp -3599
transform 1 0 29808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp -3599
transform 1 0 31004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp -3599
transform 1 0 30268 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp -3599
transform 1 0 30544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp -3599
transform -1 0 30084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp -3599
transform -1 0 29440 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp -3599
transform -1 0 28612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp -3599
transform -1 0 28244 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp -3599
transform -1 0 27968 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp -3599
transform -1 0 26772 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp -3599
transform -1 0 25944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp -3599
transform -1 0 22632 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform -1 0 21068 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform -1 0 23552 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform 1 0 23276 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform 1 0 22816 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform 1 0 21344 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform -1 0 19228 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform -1 0 19964 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp -3599
transform 1 0 21436 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp -3599
transform -1 0 17572 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp -3599
transform 1 0 18676 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp -3599
transform -1 0 16836 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp -3599
transform 1 0 15732 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp -3599
transform -1 0 15456 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp -3599
transform -1 0 18216 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp -3599
transform -1 0 19412 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp -3599
transform -1 0 20240 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp -3599
transform -1 0 17204 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp -3599
transform -1 0 16560 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp -3599
transform -1 0 16192 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp -3599
transform -1 0 22632 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp -3599
transform -1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp -3599
transform -1 0 20424 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp -3599
transform -1 0 24840 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp -3599
transform -1 0 23368 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp -3599
transform -1 0 23184 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp -3599
transform -1 0 25024 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp -3599
transform -1 0 22264 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp -3599
transform 1 0 20424 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp -3599
transform -1 0 21344 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp -3599
transform 1 0 20608 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp -3599
transform 1 0 25484 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp -3599
transform -1 0 30268 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp -3599
transform -1 0 29440 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp -3599
transform -1 0 28888 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp -3599
transform 1 0 28704 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp -3599
transform 1 0 26312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp -3599
transform -1 0 27692 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp -3599
transform -1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp -3599
transform -1 0 29624 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp -3599
transform 1 0 29624 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_42
timestamp -3599
transform -1 0 31004 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_43
timestamp -3599
transform 1 0 30084 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3
timestamp -3599
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6
timestamp -3599
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9
timestamp -3599
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12
timestamp -3599
transform 1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15
timestamp -3599
transform 1 0 2484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18
timestamp -3599
transform 1 0 2760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21
timestamp -3599
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24
timestamp -3599
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29
timestamp -3599
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp -3599
transform 1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35
timestamp -3599
transform 1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38
timestamp -3599
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41
timestamp -3599
transform 1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44
timestamp -3599
transform 1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47
timestamp -3599
transform 1 0 5428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50
timestamp -3599
transform 1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -3599
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp -3599
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60
timestamp -3599
transform 1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63
timestamp -3599
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66
timestamp -3599
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69
timestamp -3599
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72
timestamp -3599
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75
timestamp -3599
transform 1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_78
timestamp -3599
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -3599
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85
timestamp -3599
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_88
timestamp -3599
transform 1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_91
timestamp -3599
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_94
timestamp -3599
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_97
timestamp -3599
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100
timestamp -3599
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_103
timestamp -3599
transform 1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_106
timestamp -3599
transform 1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -3599
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp -3599
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_116
timestamp -3599
transform 1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119
timestamp -3599
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_122
timestamp -3599
transform 1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_125
timestamp -3599
transform 1 0 12604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_128
timestamp -3599
transform 1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_131
timestamp -3599
transform 1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_134
timestamp -3599
transform 1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp -3599
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141
timestamp -3599
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_144
timestamp -3599
transform 1 0 14352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_147
timestamp -3599
transform 1 0 14628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_150
timestamp -3599
transform 1 0 14904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_153
timestamp -3599
transform 1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156
timestamp -3599
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_159
timestamp -3599
transform 1 0 15732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_162
timestamp -3599
transform 1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -3599
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp -3599
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp -3599
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp -3599
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp -3599
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp -3599
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp -3599
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_341
timestamp -3599
transform 1 0 32476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_344
timestamp -3599
transform 1 0 32752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_347
timestamp -3599
transform 1 0 33028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_350
timestamp -3599
transform 1 0 33304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_353
timestamp -3599
transform 1 0 33580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_356
timestamp -3599
transform 1 0 33856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_359
timestamp -3599
transform 1 0 34132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp -3599
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_365
timestamp -3599
transform 1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_368
timestamp -3599
transform 1 0 34960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_371
timestamp -3599
transform 1 0 35236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_374
timestamp -3599
transform 1 0 35512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_377
timestamp -3599
transform 1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_380
timestamp -3599
transform 1 0 36064 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_383
timestamp -3599
transform 1 0 36340 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp -3599
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp -3599
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_6
timestamp -3599
transform 1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_9
timestamp -3599
transform 1 0 1932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_12
timestamp -3599
transform 1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_15
timestamp -3599
transform 1 0 2484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_18
timestamp -3599
transform 1 0 2760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_21
timestamp -3599
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_24
timestamp -3599
transform 1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_27
timestamp -3599
transform 1 0 3588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_30
timestamp -3599
transform 1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_33
timestamp -3599
transform 1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_36
timestamp -3599
transform 1 0 4416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_39
timestamp -3599
transform 1 0 4692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_42
timestamp -3599
transform 1 0 4968 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_45
timestamp -3599
transform 1 0 5244 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_48
timestamp -3599
transform 1 0 5520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_51
timestamp -3599
transform 1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp -3599
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp -3599
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_60
timestamp -3599
transform 1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_63
timestamp -3599
transform 1 0 6900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_66
timestamp -3599
transform 1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_69
timestamp -3599
transform 1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_72
timestamp -3599
transform 1 0 7728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_75
timestamp -3599
transform 1 0 8004 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_78
timestamp -3599
transform 1 0 8280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_81
timestamp -3599
transform 1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_84
timestamp -3599
transform 1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_87
timestamp -3599
transform 1 0 9108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_90
timestamp -3599
transform 1 0 9384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_93
timestamp -3599
transform 1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_96
timestamp -3599
transform 1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_99
timestamp -3599
transform 1 0 10212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_102
timestamp -3599
transform 1 0 10488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_105
timestamp -3599
transform 1 0 10764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_108
timestamp -3599
transform 1 0 11040 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp -3599
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp -3599
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_116
timestamp -3599
transform 1 0 11776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_119
timestamp -3599
transform 1 0 12052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_122
timestamp -3599
transform 1 0 12328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_125
timestamp -3599
transform 1 0 12604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_128
timestamp -3599
transform 1 0 12880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_131
timestamp -3599
transform 1 0 13156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_134
timestamp -3599
transform 1 0 13432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_137
timestamp -3599
transform 1 0 13708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_140
timestamp -3599
transform 1 0 13984 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_143
timestamp -3599
transform 1 0 14260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_146
timestamp -3599
transform 1 0 14536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_149
timestamp -3599
transform 1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_152
timestamp -3599
transform 1 0 15088 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_155
timestamp -3599
transform 1 0 15364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_158
timestamp -3599
transform 1 0 15640 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_161
timestamp -3599
transform 1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_164
timestamp -3599
transform 1 0 16192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp -3599
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_169
timestamp -3599
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_172
timestamp -3599
transform 1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_175
timestamp -3599
transform 1 0 17204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_182
timestamp -3599
transform 1 0 17848 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_185
timestamp -3599
transform 1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_188
timestamp -3599
transform 1 0 18400 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_194
timestamp -3599
transform 1 0 18952 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_197
timestamp -3599
transform 1 0 19228 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_203
timestamp -3599
transform 1 0 19780 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_206
timestamp -3599
transform 1 0 20056 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_209
timestamp -3599
transform 1 0 20332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_212
timestamp -3599
transform 1 0 20608 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_215
timestamp -3599
transform 1 0 20884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_218
timestamp -3599
transform 1 0 21160 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_221
timestamp -3599
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_225
timestamp -3599
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_228
timestamp -3599
transform 1 0 22080 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_234
timestamp -3599
transform 1 0 22632 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_239
timestamp -3599
transform 1 0 23092 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_245
timestamp -3599
transform 1 0 23644 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_251
timestamp -3599
transform 1 0 24196 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_254
timestamp -3599
transform 1 0 24472 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_257
timestamp -3599
transform 1 0 24748 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_263
timestamp -3599
transform 1 0 25300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_266
timestamp -3599
transform 1 0 25576 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_276
timestamp -3599
transform 1 0 26496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp -3599
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp -3599
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_287
timestamp -3599
transform 1 0 27508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_290
timestamp -3599
transform 1 0 27784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_293
timestamp -3599
transform 1 0 28060 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_303
timestamp -3599
transform 1 0 28980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_306
timestamp -3599
transform 1 0 29256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_311
timestamp -3599
transform 1 0 29716 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_314
timestamp -3599
transform 1 0 29992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_317
timestamp -3599
transform 1 0 30268 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_323
timestamp -3599
transform 1 0 30820 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_329
timestamp -3599
transform 1 0 31372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_332
timestamp -3599
transform 1 0 31648 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp -3599
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_337
timestamp -3599
transform 1 0 32108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_340
timestamp -3599
transform 1 0 32384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_343
timestamp -3599
transform 1 0 32660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_346
timestamp -3599
transform 1 0 32936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_349
timestamp -3599
transform 1 0 33212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_352
timestamp -3599
transform 1 0 33488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_355
timestamp -3599
transform 1 0 33764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_358
timestamp -3599
transform 1 0 34040 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_361
timestamp -3599
transform 1 0 34316 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_364
timestamp -3599
transform 1 0 34592 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_367
timestamp -3599
transform 1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_370
timestamp -3599
transform 1 0 35144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_373
timestamp -3599
transform 1 0 35420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_376
timestamp -3599
transform 1 0 35696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_379
timestamp -3599
transform 1 0 35972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_382
timestamp -3599
transform 1 0 36248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_385
timestamp -3599
transform 1 0 36524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_388
timestamp -3599
transform 1 0 36800 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp -3599
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp -3599
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp -3599
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_6
timestamp -3599
transform 1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_9
timestamp -3599
transform 1 0 1932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_12
timestamp -3599
transform 1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_15
timestamp -3599
transform 1 0 2484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_18
timestamp -3599
transform 1 0 2760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_21
timestamp -3599
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_24
timestamp -3599
transform 1 0 3312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_32
timestamp -3599
transform 1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_35
timestamp -3599
transform 1 0 4324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_38
timestamp -3599
transform 1 0 4600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_41
timestamp -3599
transform 1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_44
timestamp -3599
transform 1 0 5152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_47
timestamp -3599
transform 1 0 5428 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_50
timestamp -3599
transform 1 0 5704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_53
timestamp -3599
transform 1 0 5980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_56
timestamp -3599
transform 1 0 6256 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_59
timestamp -3599
transform 1 0 6532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_62
timestamp -3599
transform 1 0 6808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_65
timestamp -3599
transform 1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_68
timestamp -3599
transform 1 0 7360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_71
timestamp -3599
transform 1 0 7636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_74
timestamp -3599
transform 1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_77
timestamp -3599
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_80
timestamp -3599
transform 1 0 8464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp -3599
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_85
timestamp -3599
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_88
timestamp -3599
transform 1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_91
timestamp -3599
transform 1 0 9476 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_94
timestamp -3599
transform 1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_97
timestamp -3599
transform 1 0 10028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_100
timestamp -3599
transform 1 0 10304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_103
timestamp -3599
transform 1 0 10580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_106
timestamp -3599
transform 1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_109
timestamp -3599
transform 1 0 11132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_112
timestamp -3599
transform 1 0 11408 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_115
timestamp -3599
transform 1 0 11684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_118
timestamp -3599
transform 1 0 11960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_121
timestamp -3599
transform 1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_124
timestamp -3599
transform 1 0 12512 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_127
timestamp -3599
transform 1 0 12788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_130
timestamp -3599
transform 1 0 13064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_133
timestamp -3599
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_136
timestamp -3599
transform 1 0 13616 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp -3599
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_141
timestamp -3599
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_144
timestamp -3599
transform 1 0 14352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_147
timestamp -3599
transform 1 0 14628 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_150
timestamp -3599
transform 1 0 14904 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_153
timestamp -3599
transform 1 0 15180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_156
timestamp -3599
transform 1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_159
timestamp -3599
transform 1 0 15732 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_162
timestamp -3599
transform 1 0 16008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_165
timestamp -3599
transform 1 0 16284 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_169
timestamp -3599
transform 1 0 16652 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_174
timestamp -3599
transform 1 0 17112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_177
timestamp -3599
transform 1 0 17388 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_184
timestamp -3599
transform 1 0 18032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_187
timestamp -3599
transform 1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_190
timestamp -3599
transform 1 0 18584 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_193
timestamp -3599
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp -3599
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_200
timestamp -3599
transform 1 0 19504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_203
timestamp -3599
transform 1 0 19780 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_206
timestamp -3599
transform 1 0 20056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_209
timestamp -3599
transform 1 0 20332 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_212
timestamp -3599
transform 1 0 20608 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_220
timestamp -3599
transform 1 0 21344 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_226
timestamp -3599
transform 1 0 21896 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_231
timestamp -3599
transform 1 0 22356 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_237
timestamp -3599
transform 1 0 22908 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp -3599
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_260
timestamp -3599
transform 1 0 25024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_263
timestamp -3599
transform 1 0 25300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_266
timestamp -3599
transform 1 0 25576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_269
timestamp -3599
transform 1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_272
timestamp -3599
transform 1 0 26128 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_275
timestamp -3599
transform 1 0 26404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_278
timestamp -3599
transform 1 0 26680 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_281
timestamp -3599
transform 1 0 26956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_284
timestamp -3599
transform 1 0 27232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_287
timestamp -3599
transform 1 0 27508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_290
timestamp -3599
transform 1 0 27784 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_293
timestamp -3599
transform 1 0 28060 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_296
timestamp -3599
transform 1 0 28336 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_299
timestamp -3599
transform 1 0 28612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_305
timestamp -3599
transform 1 0 29164 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_317
timestamp -3599
transform 1 0 30268 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_320
timestamp -3599
transform 1 0 30544 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_323
timestamp -3599
transform 1 0 30820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_326
timestamp -3599
transform 1 0 31096 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_329
timestamp -3599
transform 1 0 31372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_332
timestamp -3599
transform 1 0 31648 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_335
timestamp -3599
transform 1 0 31924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_338
timestamp -3599
transform 1 0 32200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_341
timestamp -3599
transform 1 0 32476 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_344
timestamp -3599
transform 1 0 32752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_347
timestamp -3599
transform 1 0 33028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_350
timestamp -3599
transform 1 0 33304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_353
timestamp -3599
transform 1 0 33580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_356
timestamp -3599
transform 1 0 33856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_359
timestamp -3599
transform 1 0 34132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp -3599
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_365
timestamp -3599
transform 1 0 34684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_368
timestamp -3599
transform 1 0 34960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_371
timestamp -3599
transform 1 0 35236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_374
timestamp -3599
transform 1 0 35512 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_377
timestamp -3599
transform 1 0 35788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_380
timestamp -3599
transform 1 0 36064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_383
timestamp -3599
transform 1 0 36340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_386
timestamp -3599
transform 1 0 36616 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_389
timestamp -3599
transform 1 0 36892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_392
timestamp -3599
transform 1 0 37168 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_395
timestamp -3599
transform 1 0 37444 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_398
timestamp -3599
transform 1 0 37720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp -3599
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_6
timestamp -3599
transform 1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_9
timestamp -3599
transform 1 0 1932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_12
timestamp -3599
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_15
timestamp -3599
transform 1 0 2484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_18
timestamp -3599
transform 1 0 2760 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_22
timestamp -3599
transform 1 0 3128 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_25
timestamp -3599
transform 1 0 3404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_28
timestamp -3599
transform 1 0 3680 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_31
timestamp -3599
transform 1 0 3956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_34
timestamp -3599
transform 1 0 4232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_37
timestamp -3599
transform 1 0 4508 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_40
timestamp -3599
transform 1 0 4784 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_43
timestamp -3599
transform 1 0 5060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_46
timestamp -3599
transform 1 0 5336 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_49
timestamp -3599
transform 1 0 5612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_52
timestamp -3599
transform 1 0 5888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp -3599
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_57
timestamp -3599
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_60
timestamp -3599
transform 1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_63
timestamp -3599
transform 1 0 6900 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_66
timestamp -3599
transform 1 0 7176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_69
timestamp -3599
transform 1 0 7452 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_72
timestamp -3599
transform 1 0 7728 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_75
timestamp -3599
transform 1 0 8004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_78
timestamp -3599
transform 1 0 8280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_81
timestamp -3599
transform 1 0 8556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_84
timestamp -3599
transform 1 0 8832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_87
timestamp -3599
transform 1 0 9108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_90
timestamp -3599
transform 1 0 9384 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_93
timestamp -3599
transform 1 0 9660 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_96
timestamp -3599
transform 1 0 9936 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_99
timestamp -3599
transform 1 0 10212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_102
timestamp -3599
transform 1 0 10488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_105
timestamp -3599
transform 1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_108
timestamp -3599
transform 1 0 11040 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp -3599
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_113
timestamp -3599
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_116
timestamp -3599
transform 1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp -3599
transform 1 0 12052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_122
timestamp -3599
transform 1 0 12328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_125
timestamp -3599
transform 1 0 12604 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_128
timestamp -3599
transform 1 0 12880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_131
timestamp -3599
transform 1 0 13156 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_134
timestamp -3599
transform 1 0 13432 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_137
timestamp -3599
transform 1 0 13708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_140
timestamp -3599
transform 1 0 13984 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_143
timestamp -3599
transform 1 0 14260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_146
timestamp -3599
transform 1 0 14536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_149
timestamp -3599
transform 1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_152
timestamp -3599
transform 1 0 15088 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_155
timestamp -3599
transform 1 0 15364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_158
timestamp -3599
transform 1 0 15640 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_164
timestamp -3599
transform 1 0 16192 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp -3599
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_169
timestamp -3599
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_172
timestamp -3599
transform 1 0 16928 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_175
timestamp -3599
transform 1 0 17204 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_178
timestamp -3599
transform 1 0 17480 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_181
timestamp -3599
transform 1 0 17756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_184
timestamp -3599
transform 1 0 18032 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_187
timestamp -3599
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_190
timestamp -3599
transform 1 0 18584 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_193
timestamp -3599
transform 1 0 18860 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_200
timestamp -3599
transform 1 0 19504 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_203
timestamp -3599
transform 1 0 19780 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_206
timestamp -3599
transform 1 0 20056 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_209
timestamp -3599
transform 1 0 20332 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_212
timestamp -3599
transform 1 0 20608 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_215
timestamp -3599
transform 1 0 20884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_218
timestamp -3599
transform 1 0 21160 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_221
timestamp -3599
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_230
timestamp -3599
transform 1 0 22264 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_233
timestamp -3599
transform 1 0 22540 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_236
timestamp -3599
transform 1 0 22816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_239
timestamp -3599
transform 1 0 23092 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_242
timestamp -3599
transform 1 0 23368 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_245
timestamp -3599
transform 1 0 23644 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_248
timestamp -3599
transform 1 0 23920 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_251
timestamp -3599
transform 1 0 24196 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_254
timestamp -3599
transform 1 0 24472 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_257
timestamp -3599
transform 1 0 24748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_260
timestamp -3599
transform 1 0 25024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_263
timestamp -3599
transform 1 0 25300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_270
timestamp -3599
transform 1 0 25944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_273
timestamp -3599
transform 1 0 26220 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp -3599
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_281
timestamp -3599
transform 1 0 26956 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_285
timestamp -3599
transform 1 0 27324 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_288
timestamp -3599
transform 1 0 27600 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_292
timestamp -3599
transform 1 0 27968 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_299
timestamp -3599
transform 1 0 28612 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_328
timestamp -3599
transform 1 0 31280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_331
timestamp -3599
transform 1 0 31556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp -3599
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_337
timestamp -3599
transform 1 0 32108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_340
timestamp -3599
transform 1 0 32384 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_343
timestamp -3599
transform 1 0 32660 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_346
timestamp -3599
transform 1 0 32936 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_349
timestamp -3599
transform 1 0 33212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_352
timestamp -3599
transform 1 0 33488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_355
timestamp -3599
transform 1 0 33764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_358
timestamp -3599
transform 1 0 34040 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_361
timestamp -3599
transform 1 0 34316 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_364
timestamp -3599
transform 1 0 34592 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_367
timestamp -3599
transform 1 0 34868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_370
timestamp -3599
transform 1 0 35144 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_373
timestamp -3599
transform 1 0 35420 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_376
timestamp -3599
transform 1 0 35696 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_379
timestamp -3599
transform 1 0 35972 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_382
timestamp -3599
transform 1 0 36248 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_385
timestamp -3599
transform 1 0 36524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_388
timestamp -3599
transform 1 0 36800 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp -3599
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_393
timestamp -3599
transform 1 0 37260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_396
timestamp -3599
transform 1 0 37536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp -3599
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_6
timestamp -3599
transform 1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_9
timestamp -3599
transform 1 0 1932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_12
timestamp -3599
transform 1 0 2208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_15
timestamp -3599
transform 1 0 2484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_18
timestamp -3599
transform 1 0 2760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_21
timestamp -3599
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_24
timestamp -3599
transform 1 0 3312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -3599
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp -3599
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_32
timestamp -3599
transform 1 0 4048 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_37
timestamp -3599
transform 1 0 4508 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_40
timestamp -3599
transform 1 0 4784 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_43
timestamp -3599
transform 1 0 5060 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_46
timestamp -3599
transform 1 0 5336 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_49
timestamp -3599
transform 1 0 5612 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_52
timestamp -3599
transform 1 0 5888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_55
timestamp -3599
transform 1 0 6164 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_58
timestamp -3599
transform 1 0 6440 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_61
timestamp -3599
transform 1 0 6716 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_64
timestamp -3599
transform 1 0 6992 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_67
timestamp -3599
transform 1 0 7268 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_70
timestamp -3599
transform 1 0 7544 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_73
timestamp -3599
transform 1 0 7820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_76
timestamp -3599
transform 1 0 8096 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_79
timestamp -3599
transform 1 0 8372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp -3599
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_85
timestamp -3599
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_88
timestamp -3599
transform 1 0 9200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_91
timestamp -3599
transform 1 0 9476 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_94
timestamp -3599
transform 1 0 9752 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_97
timestamp -3599
transform 1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_100
timestamp -3599
transform 1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_103
timestamp -3599
transform 1 0 10580 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_106
timestamp -3599
transform 1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_109
timestamp -3599
transform 1 0 11132 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_112
timestamp -3599
transform 1 0 11408 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_115
timestamp -3599
transform 1 0 11684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_118
timestamp -3599
transform 1 0 11960 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_121
timestamp -3599
transform 1 0 12236 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_124
timestamp -3599
transform 1 0 12512 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_127
timestamp -3599
transform 1 0 12788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_130
timestamp -3599
transform 1 0 13064 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_133
timestamp -3599
transform 1 0 13340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_136
timestamp -3599
transform 1 0 13616 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp -3599
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_141
timestamp -3599
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_144
timestamp -3599
transform 1 0 14352 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_147
timestamp -3599
transform 1 0 14628 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_150
timestamp -3599
transform 1 0 14904 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_157
timestamp -3599
transform 1 0 15548 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_160
timestamp -3599
transform 1 0 15824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_163
timestamp -3599
transform 1 0 16100 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_166
timestamp -3599
transform 1 0 16376 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_169
timestamp -3599
transform 1 0 16652 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_172
timestamp -3599
transform 1 0 16928 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_175
timestamp -3599
transform 1 0 17204 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_178
timestamp -3599
transform 1 0 17480 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_181
timestamp -3599
transform 1 0 17756 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_184
timestamp -3599
transform 1 0 18032 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_187
timestamp -3599
transform 1 0 18308 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_190
timestamp -3599
transform 1 0 18584 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp -3599
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_202
timestamp -3599
transform 1 0 19688 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_205
timestamp -3599
transform 1 0 19964 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_208
timestamp -3599
transform 1 0 20240 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_211
timestamp -3599
transform 1 0 20516 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_214
timestamp -3599
transform 1 0 20792 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_217
timestamp -3599
transform 1 0 21068 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_225
timestamp -3599
transform 1 0 21804 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_228
timestamp -3599
transform 1 0 22080 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_231
timestamp -3599
transform 1 0 22356 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_234
timestamp -3599
transform 1 0 22632 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_237
timestamp -3599
transform 1 0 22908 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_240
timestamp -3599
transform 1 0 23184 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_247
timestamp -3599
transform 1 0 23828 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp -3599
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_253
timestamp -3599
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_256
timestamp -3599
transform 1 0 24656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_259
timestamp -3599
transform 1 0 24932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_262
timestamp -3599
transform 1 0 25208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_265
timestamp -3599
transform 1 0 25484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_268
timestamp -3599
transform 1 0 25760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_271
timestamp -3599
transform 1 0 26036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_274
timestamp -3599
transform 1 0 26312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_277
timestamp -3599
transform 1 0 26588 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_280
timestamp -3599
transform 1 0 26864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_283
timestamp -3599
transform 1 0 27140 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_286
timestamp -3599
transform 1 0 27416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_297
timestamp -3599
transform 1 0 28428 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_300
timestamp -3599
transform 1 0 28704 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_304
timestamp -3599
transform 1 0 29072 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp -3599
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_312
timestamp -3599
transform 1 0 29808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_315
timestamp -3599
transform 1 0 30084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_318
timestamp -3599
transform 1 0 30360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_321
timestamp -3599
transform 1 0 30636 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_325
timestamp -3599
transform 1 0 31004 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_328
timestamp -3599
transform 1 0 31280 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_331
timestamp -3599
transform 1 0 31556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_334
timestamp -3599
transform 1 0 31832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_337
timestamp -3599
transform 1 0 32108 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_340
timestamp -3599
transform 1 0 32384 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_343
timestamp -3599
transform 1 0 32660 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_346
timestamp -3599
transform 1 0 32936 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_349
timestamp -3599
transform 1 0 33212 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_352
timestamp -3599
transform 1 0 33488 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_355
timestamp -3599
transform 1 0 33764 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_358
timestamp -3599
transform 1 0 34040 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_361
timestamp -3599
transform 1 0 34316 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_365
timestamp -3599
transform 1 0 34684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_368
timestamp -3599
transform 1 0 34960 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_371
timestamp -3599
transform 1 0 35236 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_374
timestamp -3599
transform 1 0 35512 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_377
timestamp -3599
transform 1 0 35788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_380
timestamp -3599
transform 1 0 36064 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_383
timestamp -3599
transform 1 0 36340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_386
timestamp -3599
transform 1 0 36616 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_389
timestamp -3599
transform 1 0 36892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_392
timestamp -3599
transform 1 0 37168 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_395
timestamp -3599
transform 1 0 37444 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_398
timestamp -3599
transform 1 0 37720 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp -3599
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_6
timestamp -3599
transform 1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_9
timestamp -3599
transform 1 0 1932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_12
timestamp -3599
transform 1 0 2208 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_15
timestamp -3599
transform 1 0 2484 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_18
timestamp -3599
transform 1 0 2760 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_21
timestamp -3599
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_24
timestamp -3599
transform 1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_27
timestamp -3599
transform 1 0 3588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_30
timestamp -3599
transform 1 0 3864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_42
timestamp -3599
transform 1 0 4968 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_45
timestamp -3599
transform 1 0 5244 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_51
timestamp -3599
transform 1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp -3599
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_57
timestamp -3599
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_60
timestamp -3599
transform 1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_63
timestamp -3599
transform 1 0 6900 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_66
timestamp -3599
transform 1 0 7176 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_69
timestamp -3599
transform 1 0 7452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_72
timestamp -3599
transform 1 0 7728 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_75
timestamp -3599
transform 1 0 8004 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_78
timestamp -3599
transform 1 0 8280 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_81
timestamp -3599
transform 1 0 8556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_84
timestamp -3599
transform 1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_87
timestamp -3599
transform 1 0 9108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_90
timestamp -3599
transform 1 0 9384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_93
timestamp -3599
transform 1 0 9660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_96
timestamp -3599
transform 1 0 9936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_99
timestamp -3599
transform 1 0 10212 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_102
timestamp -3599
transform 1 0 10488 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_105
timestamp -3599
transform 1 0 10764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_108
timestamp -3599
transform 1 0 11040 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp -3599
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_113
timestamp -3599
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_116
timestamp -3599
transform 1 0 11776 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_119
timestamp -3599
transform 1 0 12052 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_122
timestamp -3599
transform 1 0 12328 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_125
timestamp -3599
transform 1 0 12604 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_128
timestamp -3599
transform 1 0 12880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_131
timestamp -3599
transform 1 0 13156 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_134
timestamp -3599
transform 1 0 13432 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_149
timestamp -3599
transform 1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_152
timestamp -3599
transform 1 0 15088 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_155
timestamp -3599
transform 1 0 15364 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_158
timestamp -3599
transform 1 0 15640 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_161
timestamp -3599
transform 1 0 15916 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_164
timestamp -3599
transform 1 0 16192 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp -3599
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_169
timestamp -3599
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_172
timestamp -3599
transform 1 0 16928 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp -3599
transform 1 0 17204 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_182
timestamp -3599
transform 1 0 17848 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_185
timestamp -3599
transform 1 0 18124 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_188
timestamp -3599
transform 1 0 18400 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_191
timestamp -3599
transform 1 0 18676 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_194
timestamp -3599
transform 1 0 18952 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_197
timestamp -3599
transform 1 0 19228 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_200
timestamp -3599
transform 1 0 19504 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_208
timestamp -3599
transform 1 0 20240 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_211
timestamp -3599
transform 1 0 20516 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_214
timestamp -3599
transform 1 0 20792 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_217
timestamp -3599
transform 1 0 21068 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_220
timestamp -3599
transform 1 0 21344 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp -3599
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp -3599
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_228
timestamp -3599
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_231
timestamp -3599
transform 1 0 22356 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_234
timestamp -3599
transform 1 0 22632 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_246
timestamp -3599
transform 1 0 23736 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_249
timestamp -3599
transform 1 0 24012 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_252
timestamp -3599
transform 1 0 24288 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_255
timestamp -3599
transform 1 0 24564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_258
timestamp -3599
transform 1 0 24840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_261
timestamp -3599
transform 1 0 25116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_264
timestamp -3599
transform 1 0 25392 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_267
timestamp -3599
transform 1 0 25668 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_270
timestamp -3599
transform 1 0 25944 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_273
timestamp -3599
transform 1 0 26220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_276
timestamp -3599
transform 1 0 26496 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp -3599
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_281
timestamp -3599
transform 1 0 26956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_284
timestamp -3599
transform 1 0 27232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_287
timestamp -3599
transform 1 0 27508 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_290
timestamp -3599
transform 1 0 27784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_293
timestamp -3599
transform 1 0 28060 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_296
timestamp -3599
transform 1 0 28336 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_299
timestamp -3599
transform 1 0 28612 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_302
timestamp -3599
transform 1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_305
timestamp -3599
transform 1 0 29164 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_308
timestamp -3599
transform 1 0 29440 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_311
timestamp -3599
transform 1 0 29716 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_314
timestamp -3599
transform 1 0 29992 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_317
timestamp -3599
transform 1 0 30268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_320
timestamp -3599
transform 1 0 30544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_323
timestamp -3599
transform 1 0 30820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_326
timestamp -3599
transform 1 0 31096 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_329
timestamp -3599
transform 1 0 31372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_332
timestamp -3599
transform 1 0 31648 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp -3599
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_337
timestamp -3599
transform 1 0 32108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_340
timestamp -3599
transform 1 0 32384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_343
timestamp -3599
transform 1 0 32660 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_348
timestamp -3599
transform 1 0 33120 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_351
timestamp -3599
transform 1 0 33396 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_354
timestamp -3599
transform 1 0 33672 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_357
timestamp -3599
transform 1 0 33948 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_360
timestamp -3599
transform 1 0 34224 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_363
timestamp -3599
transform 1 0 34500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_366
timestamp -3599
transform 1 0 34776 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_369
timestamp -3599
transform 1 0 35052 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_372
timestamp -3599
transform 1 0 35328 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_375
timestamp -3599
transform 1 0 35604 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_378
timestamp -3599
transform 1 0 35880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_381
timestamp -3599
transform 1 0 36156 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_384
timestamp -3599
transform 1 0 36432 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_387
timestamp -3599
transform 1 0 36708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_390
timestamp -3599
transform 1 0 36984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_393
timestamp -3599
transform 1 0 37260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_396
timestamp -3599
transform 1 0 37536 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp -3599
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_6
timestamp -3599
transform 1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_9
timestamp -3599
transform 1 0 1932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_12
timestamp -3599
transform 1 0 2208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_15
timestamp -3599
transform 1 0 2484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_18
timestamp -3599
transform 1 0 2760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_21
timestamp -3599
transform 1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_24
timestamp -3599
transform 1 0 3312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -3599
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_29
timestamp -3599
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_32
timestamp -3599
transform 1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_35
timestamp -3599
transform 1 0 4324 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_38
timestamp -3599
transform 1 0 4600 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_41
timestamp -3599
transform 1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_44
timestamp -3599
transform 1 0 5152 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_47
timestamp -3599
transform 1 0 5428 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_50
timestamp -3599
transform 1 0 5704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_56
timestamp -3599
transform 1 0 6256 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_59
timestamp -3599
transform 1 0 6532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_62
timestamp -3599
transform 1 0 6808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_65
timestamp -3599
transform 1 0 7084 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_70
timestamp -3599
transform 1 0 7544 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_73
timestamp -3599
transform 1 0 7820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_76
timestamp -3599
transform 1 0 8096 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_79
timestamp -3599
transform 1 0 8372 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp -3599
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_85
timestamp -3599
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_88
timestamp -3599
transform 1 0 9200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_91
timestamp -3599
transform 1 0 9476 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_94
timestamp -3599
transform 1 0 9752 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_97
timestamp -3599
transform 1 0 10028 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_100
timestamp -3599
transform 1 0 10304 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_103
timestamp -3599
transform 1 0 10580 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_106
timestamp -3599
transform 1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_109
timestamp -3599
transform 1 0 11132 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_112
timestamp -3599
transform 1 0 11408 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_115
timestamp -3599
transform 1 0 11684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_118
timestamp -3599
transform 1 0 11960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_121
timestamp -3599
transform 1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_124
timestamp -3599
transform 1 0 12512 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_134
timestamp -3599
transform 1 0 13432 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp -3599
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_144
timestamp -3599
transform 1 0 14352 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_147
timestamp -3599
transform 1 0 14628 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_150
timestamp -3599
transform 1 0 14904 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_153
timestamp -3599
transform 1 0 15180 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_156
timestamp -3599
transform 1 0 15456 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_159
timestamp -3599
transform 1 0 15732 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_162
timestamp -3599
transform 1 0 16008 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_165
timestamp -3599
transform 1 0 16284 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_168
timestamp -3599
transform 1 0 16560 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_171
timestamp -3599
transform 1 0 16836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_174
timestamp -3599
transform 1 0 17112 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_177
timestamp -3599
transform 1 0 17388 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_180
timestamp -3599
transform 1 0 17664 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_183
timestamp -3599
transform 1 0 17940 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_186
timestamp -3599
transform 1 0 18216 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_189
timestamp -3599
transform 1 0 18492 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_197
timestamp -3599
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_200
timestamp -3599
transform 1 0 19504 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_203
timestamp -3599
transform 1 0 19780 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_206
timestamp -3599
transform 1 0 20056 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_209
timestamp -3599
transform 1 0 20332 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_212
timestamp -3599
transform 1 0 20608 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_215
timestamp -3599
transform 1 0 20884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_218
timestamp -3599
transform 1 0 21160 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_226
timestamp -3599
transform 1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_229
timestamp -3599
transform 1 0 22172 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_232
timestamp -3599
transform 1 0 22448 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_235
timestamp -3599
transform 1 0 22724 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_238
timestamp -3599
transform 1 0 23000 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_241
timestamp -3599
transform 1 0 23276 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_244
timestamp -3599
transform 1 0 23552 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_247
timestamp -3599
transform 1 0 23828 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp -3599
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp -3599
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_256
timestamp -3599
transform 1 0 24656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_259
timestamp -3599
transform 1 0 24932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_262
timestamp -3599
transform 1 0 25208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_265
timestamp -3599
transform 1 0 25484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_268
timestamp -3599
transform 1 0 25760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_271
timestamp -3599
transform 1 0 26036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_274
timestamp -3599
transform 1 0 26312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_277
timestamp -3599
transform 1 0 26588 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_280
timestamp -3599
transform 1 0 26864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_283
timestamp -3599
transform 1 0 27140 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_286
timestamp -3599
transform 1 0 27416 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_289
timestamp -3599
transform 1 0 27692 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_292
timestamp -3599
transform 1 0 27968 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_297
timestamp -3599
transform 1 0 28428 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_300
timestamp -3599
transform 1 0 28704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_303
timestamp -3599
transform 1 0 28980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp -3599
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_309
timestamp -3599
transform 1 0 29532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_312
timestamp -3599
transform 1 0 29808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_315
timestamp -3599
transform 1 0 30084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_318
timestamp -3599
transform 1 0 30360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_321
timestamp -3599
transform 1 0 30636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_324
timestamp -3599
transform 1 0 30912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_327
timestamp -3599
transform 1 0 31188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_330
timestamp -3599
transform 1 0 31464 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_333
timestamp -3599
transform 1 0 31740 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_336
timestamp -3599
transform 1 0 32016 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_339
timestamp -3599
transform 1 0 32292 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_342
timestamp -3599
transform 1 0 32568 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_345
timestamp -3599
transform 1 0 32844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_348
timestamp -3599
transform 1 0 33120 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_351
timestamp -3599
transform 1 0 33396 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_354
timestamp -3599
transform 1 0 33672 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_357
timestamp -3599
transform 1 0 33948 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp -3599
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_365
timestamp -3599
transform 1 0 34684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_368
timestamp -3599
transform 1 0 34960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_371
timestamp -3599
transform 1 0 35236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_377
timestamp -3599
transform 1 0 35788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_380
timestamp -3599
transform 1 0 36064 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_383
timestamp -3599
transform 1 0 36340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_386
timestamp -3599
transform 1 0 36616 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_393
timestamp -3599
transform 1 0 37260 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_396
timestamp -3599
transform 1 0 37536 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp -3599
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_6
timestamp -3599
transform 1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_9
timestamp -3599
transform 1 0 1932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_12
timestamp -3599
transform 1 0 2208 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_15
timestamp -3599
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_18
timestamp -3599
transform 1 0 2760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_21
timestamp -3599
transform 1 0 3036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_24
timestamp -3599
transform 1 0 3312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_27
timestamp -3599
transform 1 0 3588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_30
timestamp -3599
transform 1 0 3864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_33
timestamp -3599
transform 1 0 4140 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_36
timestamp -3599
transform 1 0 4416 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_39
timestamp -3599
transform 1 0 4692 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_42
timestamp -3599
transform 1 0 4968 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_45
timestamp -3599
transform 1 0 5244 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_48
timestamp -3599
transform 1 0 5520 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_51
timestamp -3599
transform 1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp -3599
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_57
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_60
timestamp -3599
transform 1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_63
timestamp -3599
transform 1 0 6900 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_66
timestamp -3599
transform 1 0 7176 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_69
timestamp -3599
transform 1 0 7452 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_72
timestamp -3599
transform 1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_75
timestamp -3599
transform 1 0 8004 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_78
timestamp -3599
transform 1 0 8280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_81
timestamp -3599
transform 1 0 8556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_84
timestamp -3599
transform 1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_87
timestamp -3599
transform 1 0 9108 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_90
timestamp -3599
transform 1 0 9384 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_95
timestamp -3599
transform 1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_98
timestamp -3599
transform 1 0 10120 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_104
timestamp -3599
transform 1 0 10672 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp -3599
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_113
timestamp -3599
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_116
timestamp -3599
transform 1 0 11776 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_119
timestamp -3599
transform 1 0 12052 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_122
timestamp -3599
transform 1 0 12328 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_125
timestamp -3599
transform 1 0 12604 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_128
timestamp -3599
transform 1 0 12880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_131
timestamp -3599
transform 1 0 13156 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_134
timestamp -3599
transform 1 0 13432 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_137
timestamp -3599
transform 1 0 13708 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_140
timestamp -3599
transform 1 0 13984 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_143
timestamp -3599
transform 1 0 14260 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_146
timestamp -3599
transform 1 0 14536 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_149
timestamp -3599
transform 1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_152
timestamp -3599
transform 1 0 15088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_155
timestamp -3599
transform 1 0 15364 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_158
timestamp -3599
transform 1 0 15640 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_161
timestamp -3599
transform 1 0 15916 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_164
timestamp -3599
transform 1 0 16192 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp -3599
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_174
timestamp -3599
transform 1 0 17112 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_177
timestamp -3599
transform 1 0 17388 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_180
timestamp -3599
transform 1 0 17664 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_183
timestamp -3599
transform 1 0 17940 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_186
timestamp -3599
transform 1 0 18216 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_189
timestamp -3599
transform 1 0 18492 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_192
timestamp -3599
transform 1 0 18768 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_195
timestamp -3599
transform 1 0 19044 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_198
timestamp -3599
transform 1 0 19320 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_201
timestamp -3599
transform 1 0 19596 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_204
timestamp -3599
transform 1 0 19872 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_207
timestamp -3599
transform 1 0 20148 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_210
timestamp -3599
transform 1 0 20424 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_213
timestamp -3599
transform 1 0 20700 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_216
timestamp -3599
transform 1 0 20976 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_219
timestamp -3599
transform 1 0 21252 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp -3599
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp -3599
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_228
timestamp -3599
transform 1 0 22080 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_231
timestamp -3599
transform 1 0 22356 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_234
timestamp -3599
transform 1 0 22632 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_237
timestamp -3599
transform 1 0 22908 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_240
timestamp -3599
transform 1 0 23184 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_243
timestamp -3599
transform 1 0 23460 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_246
timestamp -3599
transform 1 0 23736 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_249
timestamp -3599
transform 1 0 24012 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_252
timestamp -3599
transform 1 0 24288 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_255
timestamp -3599
transform 1 0 24564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_258
timestamp -3599
transform 1 0 24840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_261
timestamp -3599
transform 1 0 25116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_264
timestamp -3599
transform 1 0 25392 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_267
timestamp -3599
transform 1 0 25668 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_270
timestamp -3599
transform 1 0 25944 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_273
timestamp -3599
transform 1 0 26220 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_276
timestamp -3599
transform 1 0 26496 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp -3599
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_281
timestamp -3599
transform 1 0 26956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_284
timestamp -3599
transform 1 0 27232 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_287
timestamp -3599
transform 1 0 27508 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_290
timestamp -3599
transform 1 0 27784 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_293
timestamp -3599
transform 1 0 28060 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_296
timestamp -3599
transform 1 0 28336 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_299
timestamp -3599
transform 1 0 28612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_302
timestamp -3599
transform 1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_305
timestamp -3599
transform 1 0 29164 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_308
timestamp -3599
transform 1 0 29440 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_311
timestamp -3599
transform 1 0 29716 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_314
timestamp -3599
transform 1 0 29992 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_317
timestamp -3599
transform 1 0 30268 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_320
timestamp -3599
transform 1 0 30544 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_323
timestamp -3599
transform 1 0 30820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_326
timestamp -3599
transform 1 0 31096 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_329
timestamp -3599
transform 1 0 31372 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_332
timestamp -3599
transform 1 0 31648 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp -3599
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_337
timestamp -3599
transform 1 0 32108 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_340
timestamp -3599
transform 1 0 32384 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_343
timestamp -3599
transform 1 0 32660 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_346
timestamp -3599
transform 1 0 32936 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_349
timestamp -3599
transform 1 0 33212 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_352
timestamp -3599
transform 1 0 33488 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_355
timestamp -3599
transform 1 0 33764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_358
timestamp -3599
transform 1 0 34040 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_361
timestamp -3599
transform 1 0 34316 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_364
timestamp -3599
transform 1 0 34592 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_367
timestamp -3599
transform 1 0 34868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_370
timestamp -3599
transform 1 0 35144 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_373
timestamp -3599
transform 1 0 35420 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_376
timestamp -3599
transform 1 0 35696 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_379
timestamp -3599
transform 1 0 35972 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_382
timestamp -3599
transform 1 0 36248 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_385
timestamp -3599
transform 1 0 36524 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_388
timestamp -3599
transform 1 0 36800 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp -3599
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_393
timestamp -3599
transform 1 0 37260 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_396
timestamp -3599
transform 1 0 37536 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_6
timestamp -3599
transform 1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_9
timestamp -3599
transform 1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_12
timestamp -3599
transform 1 0 2208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_15
timestamp -3599
transform 1 0 2484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_18
timestamp -3599
transform 1 0 2760 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_21
timestamp -3599
transform 1 0 3036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_24
timestamp -3599
transform 1 0 3312 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp -3599
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_29
timestamp -3599
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_32
timestamp -3599
transform 1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_35
timestamp -3599
transform 1 0 4324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_38
timestamp -3599
transform 1 0 4600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_41
timestamp -3599
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_44
timestamp -3599
transform 1 0 5152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_47
timestamp -3599
transform 1 0 5428 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_50
timestamp -3599
transform 1 0 5704 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_53
timestamp -3599
transform 1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_56
timestamp -3599
transform 1 0 6256 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_59
timestamp -3599
transform 1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_62
timestamp -3599
transform 1 0 6808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_65
timestamp -3599
transform 1 0 7084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_74
timestamp -3599
transform 1 0 7912 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp -3599
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_88
timestamp -3599
transform 1 0 9200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_92
timestamp -3599
transform 1 0 9568 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_98
timestamp -3599
transform 1 0 10120 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_103
timestamp -3599
transform 1 0 10580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_106
timestamp -3599
transform 1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_109
timestamp -3599
transform 1 0 11132 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_112
timestamp -3599
transform 1 0 11408 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_115
timestamp -3599
transform 1 0 11684 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_118
timestamp -3599
transform 1 0 11960 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_121
timestamp -3599
transform 1 0 12236 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_124
timestamp -3599
transform 1 0 12512 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_127
timestamp -3599
transform 1 0 12788 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_130
timestamp -3599
transform 1 0 13064 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_133
timestamp -3599
transform 1 0 13340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_136
timestamp -3599
transform 1 0 13616 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp -3599
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_141
timestamp -3599
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_144
timestamp -3599
transform 1 0 14352 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_147
timestamp -3599
transform 1 0 14628 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_150
timestamp -3599
transform 1 0 14904 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_153
timestamp -3599
transform 1 0 15180 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_156
timestamp -3599
transform 1 0 15456 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_164
timestamp -3599
transform 1 0 16192 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_167
timestamp -3599
transform 1 0 16468 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_170
timestamp -3599
transform 1 0 16744 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_173
timestamp -3599
transform 1 0 17020 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_176
timestamp -3599
transform 1 0 17296 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_179
timestamp -3599
transform 1 0 17572 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_182
timestamp -3599
transform 1 0 17848 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_185
timestamp -3599
transform 1 0 18124 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_188
timestamp -3599
transform 1 0 18400 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_191
timestamp -3599
transform 1 0 18676 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp -3599
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp -3599
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_200
timestamp -3599
transform 1 0 19504 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_203
timestamp -3599
transform 1 0 19780 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_208
timestamp -3599
transform 1 0 20240 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_211
timestamp -3599
transform 1 0 20516 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_214
timestamp -3599
transform 1 0 20792 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_217
timestamp -3599
transform 1 0 21068 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_220
timestamp -3599
transform 1 0 21344 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_223
timestamp -3599
transform 1 0 21620 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_226
timestamp -3599
transform 1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_229
timestamp -3599
transform 1 0 22172 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_232
timestamp -3599
transform 1 0 22448 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_235
timestamp -3599
transform 1 0 22724 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_238
timestamp -3599
transform 1 0 23000 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_241
timestamp -3599
transform 1 0 23276 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_244
timestamp -3599
transform 1 0 23552 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_247
timestamp -3599
transform 1 0 23828 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp -3599
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_253
timestamp -3599
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_256
timestamp -3599
transform 1 0 24656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_259
timestamp -3599
transform 1 0 24932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_262
timestamp -3599
transform 1 0 25208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_265
timestamp -3599
transform 1 0 25484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_268
timestamp -3599
transform 1 0 25760 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_271
timestamp -3599
transform 1 0 26036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_277
timestamp -3599
transform 1 0 26588 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_280
timestamp -3599
transform 1 0 26864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_283
timestamp -3599
transform 1 0 27140 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_286
timestamp -3599
transform 1 0 27416 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_289
timestamp -3599
transform 1 0 27692 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_292
timestamp -3599
transform 1 0 27968 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_295
timestamp -3599
transform 1 0 28244 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_298
timestamp -3599
transform 1 0 28520 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_301
timestamp -3599
transform 1 0 28796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_304
timestamp -3599
transform 1 0 29072 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp -3599
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_309
timestamp -3599
transform 1 0 29532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_312
timestamp -3599
transform 1 0 29808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_315
timestamp -3599
transform 1 0 30084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_318
timestamp -3599
transform 1 0 30360 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_321
timestamp -3599
transform 1 0 30636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_324
timestamp -3599
transform 1 0 30912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_327
timestamp -3599
transform 1 0 31188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_330
timestamp -3599
transform 1 0 31464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_333
timestamp -3599
transform 1 0 31740 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_336
timestamp -3599
transform 1 0 32016 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_339
timestamp -3599
transform 1 0 32292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_342
timestamp -3599
transform 1 0 32568 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_345
timestamp -3599
transform 1 0 32844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_348
timestamp -3599
transform 1 0 33120 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_351
timestamp -3599
transform 1 0 33396 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_354
timestamp -3599
transform 1 0 33672 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_357
timestamp -3599
transform 1 0 33948 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_360
timestamp -3599
transform 1 0 34224 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp -3599
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_365
timestamp -3599
transform 1 0 34684 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_368
timestamp -3599
transform 1 0 34960 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_371
timestamp -3599
transform 1 0 35236 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_374
timestamp -3599
transform 1 0 35512 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_377
timestamp -3599
transform 1 0 35788 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_380
timestamp -3599
transform 1 0 36064 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_383
timestamp -3599
transform 1 0 36340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_386
timestamp -3599
transform 1 0 36616 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_389
timestamp -3599
transform 1 0 36892 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_392
timestamp -3599
transform 1 0 37168 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_395
timestamp -3599
transform 1 0 37444 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_398
timestamp -3599
transform 1 0 37720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp -3599
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6
timestamp -3599
transform 1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_9
timestamp -3599
transform 1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_12
timestamp -3599
transform 1 0 2208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_15
timestamp -3599
transform 1 0 2484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_18
timestamp -3599
transform 1 0 2760 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_21
timestamp -3599
transform 1 0 3036 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_24
timestamp -3599
transform 1 0 3312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_27
timestamp -3599
transform 1 0 3588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_30
timestamp -3599
transform 1 0 3864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_33
timestamp -3599
transform 1 0 4140 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_36
timestamp -3599
transform 1 0 4416 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_39
timestamp -3599
transform 1 0 4692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_42
timestamp -3599
transform 1 0 4968 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_45
timestamp -3599
transform 1 0 5244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_48
timestamp -3599
transform 1 0 5520 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_51
timestamp -3599
transform 1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp -3599
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp -3599
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_60
timestamp -3599
transform 1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_63
timestamp -3599
transform 1 0 6900 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_66
timestamp -3599
transform 1 0 7176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_69
timestamp -3599
transform 1 0 7452 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_72
timestamp -3599
transform 1 0 7728 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_75
timestamp -3599
transform 1 0 8004 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_78
timestamp -3599
transform 1 0 8280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_81
timestamp -3599
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_84
timestamp -3599
transform 1 0 8832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_87
timestamp -3599
transform 1 0 9108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_90
timestamp -3599
transform 1 0 9384 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_93
timestamp -3599
transform 1 0 9660 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_96
timestamp -3599
transform 1 0 9936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_99
timestamp -3599
transform 1 0 10212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_102
timestamp -3599
transform 1 0 10488 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_105
timestamp -3599
transform 1 0 10764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_108
timestamp -3599
transform 1 0 11040 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp -3599
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_113
timestamp -3599
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_116
timestamp -3599
transform 1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_119
timestamp -3599
transform 1 0 12052 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_122
timestamp -3599
transform 1 0 12328 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_125
timestamp -3599
transform 1 0 12604 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_128
timestamp -3599
transform 1 0 12880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_131
timestamp -3599
transform 1 0 13156 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_134
timestamp -3599
transform 1 0 13432 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_137
timestamp -3599
transform 1 0 13708 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_140
timestamp -3599
transform 1 0 13984 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_143
timestamp -3599
transform 1 0 14260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_146
timestamp -3599
transform 1 0 14536 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_149
timestamp -3599
transform 1 0 14812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_152
timestamp -3599
transform 1 0 15088 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_172
timestamp -3599
transform 1 0 16928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_189
timestamp -3599
transform 1 0 18492 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_193
timestamp -3599
transform 1 0 18860 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_199
timestamp -3599
transform 1 0 19412 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_214
timestamp -3599
transform 1 0 20792 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_217
timestamp -3599
transform 1 0 21068 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp -3599
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_228
timestamp -3599
transform 1 0 22080 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_234
timestamp -3599
transform 1 0 22632 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_237
timestamp -3599
transform 1 0 22908 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_240
timestamp -3599
transform 1 0 23184 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_243
timestamp -3599
transform 1 0 23460 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_248
timestamp -3599
transform 1 0 23920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_251
timestamp -3599
transform 1 0 24196 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_254
timestamp -3599
transform 1 0 24472 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_257
timestamp -3599
transform 1 0 24748 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_260
timestamp -3599
transform 1 0 25024 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_265
timestamp -3599
transform 1 0 25484 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_269
timestamp -3599
transform 1 0 25852 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp -3599
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_281
timestamp -3599
transform 1 0 26956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_284
timestamp -3599
transform 1 0 27232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_287
timestamp -3599
transform 1 0 27508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_290
timestamp -3599
transform 1 0 27784 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_293
timestamp -3599
transform 1 0 28060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_296
timestamp -3599
transform 1 0 28336 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_299
timestamp -3599
transform 1 0 28612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_302
timestamp -3599
transform 1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_305
timestamp -3599
transform 1 0 29164 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_308
timestamp -3599
transform 1 0 29440 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_311
timestamp -3599
transform 1 0 29716 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_314
timestamp -3599
transform 1 0 29992 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_317
timestamp -3599
transform 1 0 30268 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_320
timestamp -3599
transform 1 0 30544 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_323
timestamp -3599
transform 1 0 30820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_326
timestamp -3599
transform 1 0 31096 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_329
timestamp -3599
transform 1 0 31372 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_332
timestamp -3599
transform 1 0 31648 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp -3599
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_337
timestamp -3599
transform 1 0 32108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_340
timestamp -3599
transform 1 0 32384 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_343
timestamp -3599
transform 1 0 32660 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_346
timestamp -3599
transform 1 0 32936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_349
timestamp -3599
transform 1 0 33212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_352
timestamp -3599
transform 1 0 33488 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_355
timestamp -3599
transform 1 0 33764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_358
timestamp -3599
transform 1 0 34040 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_361
timestamp -3599
transform 1 0 34316 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_364
timestamp -3599
transform 1 0 34592 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_367
timestamp -3599
transform 1 0 34868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_370
timestamp -3599
transform 1 0 35144 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_373
timestamp -3599
transform 1 0 35420 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_376
timestamp -3599
transform 1 0 35696 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_379
timestamp -3599
transform 1 0 35972 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_382
timestamp -3599
transform 1 0 36248 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_385
timestamp -3599
transform 1 0 36524 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_388
timestamp -3599
transform 1 0 36800 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp -3599
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_393
timestamp -3599
transform 1 0 37260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_396
timestamp -3599
transform 1 0 37536 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_6
timestamp -3599
transform 1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_9
timestamp -3599
transform 1 0 1932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_12
timestamp -3599
transform 1 0 2208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_15
timestamp -3599
transform 1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_18
timestamp -3599
transform 1 0 2760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_21
timestamp -3599
transform 1 0 3036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_24
timestamp -3599
transform 1 0 3312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp -3599
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_32
timestamp -3599
transform 1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_35
timestamp -3599
transform 1 0 4324 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_38
timestamp -3599
transform 1 0 4600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_41
timestamp -3599
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_44
timestamp -3599
transform 1 0 5152 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_47
timestamp -3599
transform 1 0 5428 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_50
timestamp -3599
transform 1 0 5704 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_53
timestamp -3599
transform 1 0 5980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_56
timestamp -3599
transform 1 0 6256 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_59
timestamp -3599
transform 1 0 6532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_62
timestamp -3599
transform 1 0 6808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_65
timestamp -3599
transform 1 0 7084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_68
timestamp -3599
transform 1 0 7360 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_71
timestamp -3599
transform 1 0 7636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_74
timestamp -3599
transform 1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_77
timestamp -3599
transform 1 0 8188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_80
timestamp -3599
transform 1 0 8464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp -3599
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_85
timestamp -3599
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_88
timestamp -3599
transform 1 0 9200 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_91
timestamp -3599
transform 1 0 9476 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_94
timestamp -3599
transform 1 0 9752 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_97
timestamp -3599
transform 1 0 10028 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_100
timestamp -3599
transform 1 0 10304 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_103
timestamp -3599
transform 1 0 10580 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_106
timestamp -3599
transform 1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_109
timestamp -3599
transform 1 0 11132 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_112
timestamp -3599
transform 1 0 11408 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_115
timestamp -3599
transform 1 0 11684 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_118
timestamp -3599
transform 1 0 11960 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_121
timestamp -3599
transform 1 0 12236 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_124
timestamp -3599
transform 1 0 12512 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_127
timestamp -3599
transform 1 0 12788 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_130
timestamp -3599
transform 1 0 13064 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_133
timestamp -3599
transform 1 0 13340 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_136
timestamp -3599
transform 1 0 13616 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp -3599
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_141
timestamp -3599
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_144
timestamp -3599
transform 1 0 14352 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_147
timestamp -3599
transform 1 0 14628 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_150
timestamp -3599
transform 1 0 14904 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_153
timestamp -3599
transform 1 0 15180 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_156
timestamp -3599
transform 1 0 15456 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_159
timestamp -3599
transform 1 0 15732 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_162
timestamp -3599
transform 1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_165
timestamp -3599
transform 1 0 16284 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_168
timestamp -3599
transform 1 0 16560 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_171
timestamp -3599
transform 1 0 16836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_174
timestamp -3599
transform 1 0 17112 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_177
timestamp -3599
transform 1 0 17388 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_180
timestamp -3599
transform 1 0 17664 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_183
timestamp -3599
transform 1 0 17940 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_186
timestamp -3599
transform 1 0 18216 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_189
timestamp -3599
transform 1 0 18492 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_192
timestamp -3599
transform 1 0 18768 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp -3599
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_197
timestamp -3599
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_200
timestamp -3599
transform 1 0 19504 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_203
timestamp -3599
transform 1 0 19780 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_206
timestamp -3599
transform 1 0 20056 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_209
timestamp -3599
transform 1 0 20332 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_212
timestamp -3599
transform 1 0 20608 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_215
timestamp -3599
transform 1 0 20884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_218
timestamp -3599
transform 1 0 21160 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_221
timestamp -3599
transform 1 0 21436 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_224
timestamp -3599
transform 1 0 21712 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_227
timestamp -3599
transform 1 0 21988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_230
timestamp -3599
transform 1 0 22264 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_233
timestamp -3599
transform 1 0 22540 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_236
timestamp -3599
transform 1 0 22816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_239
timestamp -3599
transform 1 0 23092 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_242
timestamp -3599
transform 1 0 23368 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_245
timestamp -3599
transform 1 0 23644 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_248
timestamp -3599
transform 1 0 23920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp -3599
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_253
timestamp -3599
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_256
timestamp -3599
transform 1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_259
timestamp -3599
transform 1 0 24932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_262
timestamp -3599
transform 1 0 25208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_265
timestamp -3599
transform 1 0 25484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_268
timestamp -3599
transform 1 0 25760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_271
timestamp -3599
transform 1 0 26036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_274
timestamp -3599
transform 1 0 26312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_277
timestamp -3599
transform 1 0 26588 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_280
timestamp -3599
transform 1 0 26864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_283
timestamp -3599
transform 1 0 27140 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_286
timestamp -3599
transform 1 0 27416 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_289
timestamp -3599
transform 1 0 27692 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_292
timestamp -3599
transform 1 0 27968 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_295
timestamp -3599
transform 1 0 28244 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_298
timestamp -3599
transform 1 0 28520 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_301
timestamp -3599
transform 1 0 28796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_304
timestamp -3599
transform 1 0 29072 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp -3599
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_309
timestamp -3599
transform 1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_312
timestamp -3599
transform 1 0 29808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_315
timestamp -3599
transform 1 0 30084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_318
timestamp -3599
transform 1 0 30360 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_321
timestamp -3599
transform 1 0 30636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_324
timestamp -3599
transform 1 0 30912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_327
timestamp -3599
transform 1 0 31188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_330
timestamp -3599
transform 1 0 31464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_333
timestamp -3599
transform 1 0 31740 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_336
timestamp -3599
transform 1 0 32016 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_339
timestamp -3599
transform 1 0 32292 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_342
timestamp -3599
transform 1 0 32568 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_345
timestamp -3599
transform 1 0 32844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_348
timestamp -3599
transform 1 0 33120 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_351
timestamp -3599
transform 1 0 33396 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_354
timestamp -3599
transform 1 0 33672 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_357
timestamp -3599
transform 1 0 33948 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_360
timestamp -3599
transform 1 0 34224 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp -3599
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_365
timestamp -3599
transform 1 0 34684 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_368
timestamp -3599
transform 1 0 34960 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_371
timestamp -3599
transform 1 0 35236 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_374
timestamp -3599
transform 1 0 35512 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_377
timestamp -3599
transform 1 0 35788 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_380
timestamp -3599
transform 1 0 36064 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_383
timestamp -3599
transform 1 0 36340 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_386
timestamp -3599
transform 1 0 36616 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp -3599
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_8
timestamp -3599
transform 1 0 1840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_11
timestamp -3599
transform 1 0 2116 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_14
timestamp -3599
transform 1 0 2392 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_17
timestamp -3599
transform 1 0 2668 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_20
timestamp -3599
transform 1 0 2944 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_23
timestamp -3599
transform 1 0 3220 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_26
timestamp -3599
transform 1 0 3496 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_33
timestamp -3599
transform 1 0 4140 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_36
timestamp -3599
transform 1 0 4416 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_39
timestamp -3599
transform 1 0 4692 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_42
timestamp -3599
transform 1 0 4968 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_49
timestamp -3599
transform 1 0 5612 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_52
timestamp -3599
transform 1 0 5888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp -3599
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp -3599
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_60
timestamp -3599
transform 1 0 6624 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_63
timestamp -3599
transform 1 0 6900 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_69
timestamp -3599
transform 1 0 7452 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_72
timestamp -3599
transform 1 0 7728 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_75
timestamp -3599
transform 1 0 8004 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_78
timestamp -3599
transform 1 0 8280 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_81
timestamp -3599
transform 1 0 8556 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_89
timestamp -3599
transform 1 0 9292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_92
timestamp -3599
transform 1 0 9568 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_95
timestamp -3599
transform 1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_98
timestamp -3599
transform 1 0 10120 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_101
timestamp -3599
transform 1 0 10396 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_104
timestamp -3599
transform 1 0 10672 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_109
timestamp -3599
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp -3599
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_116
timestamp -3599
transform 1 0 11776 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_119
timestamp -3599
transform 1 0 12052 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_122
timestamp -3599
transform 1 0 12328 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_129
timestamp -3599
transform 1 0 12972 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_132
timestamp -3599
transform 1 0 13248 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_135
timestamp -3599
transform 1 0 13524 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_138
timestamp -3599
transform 1 0 13800 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_141
timestamp -3599
transform 1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_144
timestamp -3599
transform 1 0 14352 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_149
timestamp -3599
transform 1 0 14812 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_152
timestamp -3599
transform 1 0 15088 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_155
timestamp -3599
transform 1 0 15364 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_158
timestamp -3599
transform 1 0 15640 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_161
timestamp -3599
transform 1 0 15916 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_164
timestamp -3599
transform 1 0 16192 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp -3599
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_173
timestamp -3599
transform 1 0 17020 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_176
timestamp -3599
transform 1 0 17296 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_179
timestamp -3599
transform 1 0 17572 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_182
timestamp -3599
transform 1 0 17848 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_189
timestamp -3599
transform 1 0 18492 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_192
timestamp -3599
transform 1 0 18768 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_195
timestamp -3599
transform 1 0 19044 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_197
timestamp -3599
transform 1 0 19228 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_200
timestamp -3599
transform 1 0 19504 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_203
timestamp -3599
transform 1 0 19780 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_209
timestamp -3599
transform 1 0 20332 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_212
timestamp -3599
transform 1 0 20608 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_215
timestamp -3599
transform 1 0 20884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_218
timestamp -3599
transform 1 0 21160 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp -3599
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_229
timestamp -3599
transform 1 0 22172 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_232
timestamp -3599
transform 1 0 22448 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_235
timestamp -3599
transform 1 0 22724 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_238
timestamp -3599
transform 1 0 23000 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_241
timestamp -3599
transform 1 0 23276 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_244
timestamp -3599
transform 1 0 23552 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_249
timestamp -3599
transform 1 0 24012 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_253
timestamp -3599
transform 1 0 24380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_256
timestamp -3599
transform 1 0 24656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_259
timestamp -3599
transform 1 0 24932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_262
timestamp -3599
transform 1 0 25208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_269
timestamp -3599
transform 1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_272
timestamp -3599
transform 1 0 26128 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_275
timestamp -3599
transform 1 0 26404 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp -3599
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_281
timestamp -3599
transform 1 0 26956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_284
timestamp -3599
transform 1 0 27232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_289
timestamp -3599
transform 1 0 27692 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_292
timestamp -3599
transform 1 0 27968 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_295
timestamp -3599
transform 1 0 28244 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_298
timestamp -3599
transform 1 0 28520 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_301
timestamp -3599
transform 1 0 28796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_304
timestamp -3599
transform 1 0 29072 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_307
timestamp -3599
transform 1 0 29348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_313
timestamp -3599
transform 1 0 29900 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_316
timestamp -3599
transform 1 0 30176 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_319
timestamp -3599
transform 1 0 30452 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_322
timestamp -3599
transform 1 0 30728 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_329
timestamp -3599
transform 1 0 31372 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_332
timestamp -3599
transform 1 0 31648 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp -3599
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_337
timestamp -3599
transform 1 0 32108 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_340
timestamp -3599
transform 1 0 32384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_343
timestamp -3599
transform 1 0 32660 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_349
timestamp -3599
transform 1 0 33212 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_352
timestamp -3599
transform 1 0 33488 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_355
timestamp -3599
transform 1 0 33764 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_358
timestamp -3599
transform 1 0 34040 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_361
timestamp -3599
transform 1 0 34316 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_369
timestamp -3599
transform 1 0 35052 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_372
timestamp -3599
transform 1 0 35328 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_375
timestamp -3599
transform 1 0 35604 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_378
timestamp -3599
transform 1 0 35880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_389
timestamp -3599
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp -3599
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output1
timestamp -3599
transform 1 0 37444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp -3599
transform 1 0 37812 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp -3599
transform 1 0 38180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp -3599
transform 1 0 37812 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp -3599
transform 1 0 38180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp -3599
transform 1 0 37812 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp -3599
transform 1 0 38180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp -3599
transform 1 0 37812 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp -3599
transform 1 0 38180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp -3599
transform 1 0 37812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp -3599
transform 1 0 38180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp -3599
transform 1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp -3599
transform 1 0 37812 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp -3599
transform 1 0 38180 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp -3599
transform 1 0 38180 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp -3599
transform 1 0 37812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp -3599
transform 1 0 38180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp -3599
transform 1 0 37812 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp -3599
transform 1 0 37444 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp -3599
transform 1 0 37444 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp -3599
transform 1 0 37812 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp -3599
transform 1 0 37076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp -3599
transform 1 0 37444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp -3599
transform 1 0 36708 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp -3599
transform 1 0 36156 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp -3599
transform 1 0 36432 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp -3599
transform 1 0 37812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp -3599
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp -3599
transform 1 0 37812 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp -3599
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp -3599
transform 1 0 37812 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp -3599
transform 1 0 38180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp -3599
transform -1 0 4140 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp -3599
transform -1 0 22172 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp -3599
transform -1 0 24012 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp -3599
transform -1 0 25852 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp -3599
transform -1 0 27692 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp -3599
transform -1 0 29900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp -3599
transform -1 0 31372 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp -3599
transform -1 0 33212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp -3599
transform -1 0 35052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp -3599
transform -1 0 36892 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp -3599
transform 1 0 38180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp -3599
transform -1 0 5612 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp -3599
transform -1 0 7452 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp -3599
transform -1 0 9292 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp -3599
transform -1 0 11132 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp -3599
transform -1 0 12972 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp -3599
transform -1 0 14812 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp -3599
transform -1 0 17020 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp -3599
transform -1 0 18492 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp -3599
transform -1 0 20332 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp -3599
transform 1 0 16928 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp -3599
transform 1 0 17480 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp -3599
transform 1 0 17296 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp -3599
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp -3599
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp -3599
transform 1 0 18584 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp -3599
transform 1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp -3599
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp -3599
transform 1 0 19412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp -3599
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp -3599
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp -3599
transform 1 0 19964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp -3599
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp -3599
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp -3599
transform 1 0 21068 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp -3599
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp -3599
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp -3599
transform 1 0 22540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp -3599
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp -3599
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp -3599
transform 1 0 22724 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp -3599
transform 1 0 26220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp -3599
transform 1 0 25760 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp -3599
transform 1 0 26128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp -3599
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp -3599
transform 1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp -3599
transform 1 0 27692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp -3599
transform 1 0 23644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp -3599
transform 1 0 23276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp -3599
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp -3599
transform 1 0 23828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp -3599
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp -3599
transform 1 0 25116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp -3599
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp -3599
transform 1 0 24932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp -3599
transform -1 0 27508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp -3599
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp -3599
transform 1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp -3599
transform 1 0 30452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp -3599
transform 1 0 31372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp -3599
transform 1 0 31004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp -3599
transform 1 0 32108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp -3599
transform 1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp -3599
transform -1 0 28796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp -3599
transform -1 0 29164 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp -3599
transform -1 0 28612 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp -3599
transform -1 0 28980 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp -3599
transform -1 0 29900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp -3599
transform -1 0 30268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp -3599
transform -1 0 29716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp -3599
transform 1 0 30268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output105
timestamp -3599
transform -1 0 1840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp -3599
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp -3599
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp -3599
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp -3599
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_38
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_39
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_40
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_41
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_42
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_43
timestamp -3599
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_44
timestamp -3599
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_45
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_46
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_47
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_48
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_49
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_50
timestamp -3599
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_51
timestamp -3599
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_52
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_53
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_54
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_55
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_56
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_57
timestamp -3599
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_58
timestamp -3599
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_59
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_60
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_61
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_62
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_63
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_64
timestamp -3599
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_65
timestamp -3599
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_66
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_67
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_68
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_69
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_70
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_71
timestamp -3599
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_72
timestamp -3599
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_73
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_74
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_75
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_76
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_77
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_78
timestamp -3599
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp -3599
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_80
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_81
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_83
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_84
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_85
timestamp -3599
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_86
timestamp -3599
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_87
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_88
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_89
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_90
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_91
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_92
timestamp -3599
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_93
timestamp -3599
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_94
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_95
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_96
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_97
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_98
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_99
timestamp -3599
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_100
timestamp -3599
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_101
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_102
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_103
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_104
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_105
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_106
timestamp -3599
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_107
timestamp -3599
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_108
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_109
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_110
timestamp -3599
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_111
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_112
timestamp -3599
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_113
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_114
timestamp -3599
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_115
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_116
timestamp -3599
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_117
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_118
timestamp -3599
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_119
timestamp -3599
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_120
timestamp -3599
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_121
timestamp -3599
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 1096 120 1216 0 FreeSans 480 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 3816 120 3936 0 FreeSans 480 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal3 s 0 4360 120 4480 0 FreeSans 480 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal3 s 0 4632 120 4752 0 FreeSans 480 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal3 s 0 4904 120 5024 0 FreeSans 480 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal3 s 0 5176 120 5296 0 FreeSans 480 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal3 s 0 5448 120 5568 0 FreeSans 480 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal3 s 0 5720 120 5840 0 FreeSans 480 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal3 s 0 5992 120 6112 0 FreeSans 480 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal3 s 0 6264 120 6384 0 FreeSans 480 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal3 s 0 1368 120 1488 0 FreeSans 480 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal3 s 0 6536 120 6656 0 FreeSans 480 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal3 s 0 6808 120 6928 0 FreeSans 480 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal3 s 0 7080 120 7200 0 FreeSans 480 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal3 s 0 7352 120 7472 0 FreeSans 480 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal3 s 0 7624 120 7744 0 FreeSans 480 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal3 s 0 7896 120 8016 0 FreeSans 480 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal3 s 0 8440 120 8560 0 FreeSans 480 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal3 s 0 8712 120 8832 0 FreeSans 480 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal3 s 0 8984 120 9104 0 FreeSans 480 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal3 s 0 1640 120 1760 0 FreeSans 480 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal3 s 0 9256 120 9376 0 FreeSans 480 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal3 s 0 9528 120 9648 0 FreeSans 480 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal3 s 0 1912 120 2032 0 FreeSans 480 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal3 s 0 2184 120 2304 0 FreeSans 480 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal3 s 0 2456 120 2576 0 FreeSans 480 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal3 s 0 2728 120 2848 0 FreeSans 480 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal3 s 0 3000 120 3120 0 FreeSans 480 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal3 s 0 3272 120 3392 0 FreeSans 480 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal3 s 0 3544 120 3664 0 FreeSans 480 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal3 s 39808 1096 39928 1216 0 FreeSans 480 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal3 s 39808 3816 39928 3936 0 FreeSans 480 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal3 s 39808 4088 39928 4208 0 FreeSans 480 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal3 s 39808 4360 39928 4480 0 FreeSans 480 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal3 s 39808 4632 39928 4752 0 FreeSans 480 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal3 s 39808 4904 39928 5024 0 FreeSans 480 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal3 s 39808 5176 39928 5296 0 FreeSans 480 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal3 s 39808 5448 39928 5568 0 FreeSans 480 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal3 s 39808 5720 39928 5840 0 FreeSans 480 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal3 s 39808 5992 39928 6112 0 FreeSans 480 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal3 s 39808 6264 39928 6384 0 FreeSans 480 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal3 s 39808 1368 39928 1488 0 FreeSans 480 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal3 s 39808 6536 39928 6656 0 FreeSans 480 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal3 s 39808 6808 39928 6928 0 FreeSans 480 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal3 s 39808 7080 39928 7200 0 FreeSans 480 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal3 s 39808 7352 39928 7472 0 FreeSans 480 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal3 s 39808 7624 39928 7744 0 FreeSans 480 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal3 s 39808 7896 39928 8016 0 FreeSans 480 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal3 s 39808 8168 39928 8288 0 FreeSans 480 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal3 s 39808 8440 39928 8560 0 FreeSans 480 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal3 s 39808 8712 39928 8832 0 FreeSans 480 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal3 s 39808 8984 39928 9104 0 FreeSans 480 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal3 s 39808 1640 39928 1760 0 FreeSans 480 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal3 s 39808 9256 39928 9376 0 FreeSans 480 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal3 s 39808 9528 39928 9648 0 FreeSans 480 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal3 s 39808 1912 39928 2032 0 FreeSans 480 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal3 s 39808 2184 39928 2304 0 FreeSans 480 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal3 s 39808 2456 39928 2576 0 FreeSans 480 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal3 s 39808 2728 39928 2848 0 FreeSans 480 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal3 s 39808 3000 39928 3120 0 FreeSans 480 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal3 s 39808 3272 39928 3392 0 FreeSans 480 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal3 s 39808 3544 39928 3664 0 FreeSans 480 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal2 s 31758 0 31814 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal2 s 34518 0 34574 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal2 s 34794 0 34850 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal2 s 35070 0 35126 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal2 s 35346 0 35402 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal2 s 35622 0 35678 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal2 s 35898 0 35954 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal2 s 36174 0 36230 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal2 s 36450 0 36506 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal2 s 36726 0 36782 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal2 s 37002 0 37058 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal2 s 32034 0 32090 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal2 s 32310 0 32366 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal2 s 32586 0 32642 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal2 s 32862 0 32918 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal2 s 33138 0 33194 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal2 s 33414 0 33470 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal2 s 33690 0 33746 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal2 s 33966 0 34022 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal2 s 34242 0 34298 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal2 s 3330 11096 3386 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal2 s 21730 11096 21786 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal2 s 23570 11096 23626 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal2 s 25410 11096 25466 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal2 s 27250 11096 27306 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal2 s 29090 11096 29146 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal2 s 30930 11096 30986 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal2 s 32770 11096 32826 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal2 s 34610 11096 34666 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal2 s 36450 11096 36506 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal2 s 38290 11096 38346 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal2 s 5170 11096 5226 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal2 s 7010 11096 7066 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal2 s 8850 11096 8906 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal2 s 10690 11096 10746 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal2 s 12530 11096 12586 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal2 s 14370 11096 14426 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal2 s 16210 11096 16266 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal2 s 18050 11096 18106 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal2 s 19890 11096 19946 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal2 s 2778 0 2834 56 0 FreeSans 224 0 0 0 N1END[0]
port 104 nsew signal input
flabel metal2 s 3054 0 3110 56 0 FreeSans 224 0 0 0 N1END[1]
port 105 nsew signal input
flabel metal2 s 3330 0 3386 56 0 FreeSans 224 0 0 0 N1END[2]
port 106 nsew signal input
flabel metal2 s 3606 0 3662 56 0 FreeSans 224 0 0 0 N1END[3]
port 107 nsew signal input
flabel metal2 s 6090 0 6146 56 0 FreeSans 224 0 0 0 N2END[0]
port 108 nsew signal input
flabel metal2 s 6366 0 6422 56 0 FreeSans 224 0 0 0 N2END[1]
port 109 nsew signal input
flabel metal2 s 6642 0 6698 56 0 FreeSans 224 0 0 0 N2END[2]
port 110 nsew signal input
flabel metal2 s 6918 0 6974 56 0 FreeSans 224 0 0 0 N2END[3]
port 111 nsew signal input
flabel metal2 s 7194 0 7250 56 0 FreeSans 224 0 0 0 N2END[4]
port 112 nsew signal input
flabel metal2 s 7470 0 7526 56 0 FreeSans 224 0 0 0 N2END[5]
port 113 nsew signal input
flabel metal2 s 7746 0 7802 56 0 FreeSans 224 0 0 0 N2END[6]
port 114 nsew signal input
flabel metal2 s 8022 0 8078 56 0 FreeSans 224 0 0 0 N2END[7]
port 115 nsew signal input
flabel metal2 s 3882 0 3938 56 0 FreeSans 224 0 0 0 N2MID[0]
port 116 nsew signal input
flabel metal2 s 4158 0 4214 56 0 FreeSans 224 0 0 0 N2MID[1]
port 117 nsew signal input
flabel metal2 s 4434 0 4490 56 0 FreeSans 224 0 0 0 N2MID[2]
port 118 nsew signal input
flabel metal2 s 4710 0 4766 56 0 FreeSans 224 0 0 0 N2MID[3]
port 119 nsew signal input
flabel metal2 s 4986 0 5042 56 0 FreeSans 224 0 0 0 N2MID[4]
port 120 nsew signal input
flabel metal2 s 5262 0 5318 56 0 FreeSans 224 0 0 0 N2MID[5]
port 121 nsew signal input
flabel metal2 s 5538 0 5594 56 0 FreeSans 224 0 0 0 N2MID[6]
port 122 nsew signal input
flabel metal2 s 5814 0 5870 56 0 FreeSans 224 0 0 0 N2MID[7]
port 123 nsew signal input
flabel metal2 s 8298 0 8354 56 0 FreeSans 224 0 0 0 N4END[0]
port 124 nsew signal input
flabel metal2 s 11058 0 11114 56 0 FreeSans 224 0 0 0 N4END[10]
port 125 nsew signal input
flabel metal2 s 11334 0 11390 56 0 FreeSans 224 0 0 0 N4END[11]
port 126 nsew signal input
flabel metal2 s 11610 0 11666 56 0 FreeSans 224 0 0 0 N4END[12]
port 127 nsew signal input
flabel metal2 s 11886 0 11942 56 0 FreeSans 224 0 0 0 N4END[13]
port 128 nsew signal input
flabel metal2 s 12162 0 12218 56 0 FreeSans 224 0 0 0 N4END[14]
port 129 nsew signal input
flabel metal2 s 12438 0 12494 56 0 FreeSans 224 0 0 0 N4END[15]
port 130 nsew signal input
flabel metal2 s 8574 0 8630 56 0 FreeSans 224 0 0 0 N4END[1]
port 131 nsew signal input
flabel metal2 s 8850 0 8906 56 0 FreeSans 224 0 0 0 N4END[2]
port 132 nsew signal input
flabel metal2 s 9126 0 9182 56 0 FreeSans 224 0 0 0 N4END[3]
port 133 nsew signal input
flabel metal2 s 9402 0 9458 56 0 FreeSans 224 0 0 0 N4END[4]
port 134 nsew signal input
flabel metal2 s 9678 0 9734 56 0 FreeSans 224 0 0 0 N4END[5]
port 135 nsew signal input
flabel metal2 s 9954 0 10010 56 0 FreeSans 224 0 0 0 N4END[6]
port 136 nsew signal input
flabel metal2 s 10230 0 10286 56 0 FreeSans 224 0 0 0 N4END[7]
port 137 nsew signal input
flabel metal2 s 10506 0 10562 56 0 FreeSans 224 0 0 0 N4END[8]
port 138 nsew signal input
flabel metal2 s 10782 0 10838 56 0 FreeSans 224 0 0 0 N4END[9]
port 139 nsew signal input
flabel metal2 s 12714 0 12770 56 0 FreeSans 224 0 0 0 NN4END[0]
port 140 nsew signal input
flabel metal2 s 15474 0 15530 56 0 FreeSans 224 0 0 0 NN4END[10]
port 141 nsew signal input
flabel metal2 s 15750 0 15806 56 0 FreeSans 224 0 0 0 NN4END[11]
port 142 nsew signal input
flabel metal2 s 16026 0 16082 56 0 FreeSans 224 0 0 0 NN4END[12]
port 143 nsew signal input
flabel metal2 s 16302 0 16358 56 0 FreeSans 224 0 0 0 NN4END[13]
port 144 nsew signal input
flabel metal2 s 16578 0 16634 56 0 FreeSans 224 0 0 0 NN4END[14]
port 145 nsew signal input
flabel metal2 s 16854 0 16910 56 0 FreeSans 224 0 0 0 NN4END[15]
port 146 nsew signal input
flabel metal2 s 12990 0 13046 56 0 FreeSans 224 0 0 0 NN4END[1]
port 147 nsew signal input
flabel metal2 s 13266 0 13322 56 0 FreeSans 224 0 0 0 NN4END[2]
port 148 nsew signal input
flabel metal2 s 13542 0 13598 56 0 FreeSans 224 0 0 0 NN4END[3]
port 149 nsew signal input
flabel metal2 s 13818 0 13874 56 0 FreeSans 224 0 0 0 NN4END[4]
port 150 nsew signal input
flabel metal2 s 14094 0 14150 56 0 FreeSans 224 0 0 0 NN4END[5]
port 151 nsew signal input
flabel metal2 s 14370 0 14426 56 0 FreeSans 224 0 0 0 NN4END[6]
port 152 nsew signal input
flabel metal2 s 14646 0 14702 56 0 FreeSans 224 0 0 0 NN4END[7]
port 153 nsew signal input
flabel metal2 s 14922 0 14978 56 0 FreeSans 224 0 0 0 NN4END[8]
port 154 nsew signal input
flabel metal2 s 15198 0 15254 56 0 FreeSans 224 0 0 0 NN4END[9]
port 155 nsew signal input
flabel metal2 s 17130 0 17186 56 0 FreeSans 224 0 0 0 S1BEG[0]
port 156 nsew signal output
flabel metal2 s 17406 0 17462 56 0 FreeSans 224 0 0 0 S1BEG[1]
port 157 nsew signal output
flabel metal2 s 17682 0 17738 56 0 FreeSans 224 0 0 0 S1BEG[2]
port 158 nsew signal output
flabel metal2 s 17958 0 18014 56 0 FreeSans 224 0 0 0 S1BEG[3]
port 159 nsew signal output
flabel metal2 s 18234 0 18290 56 0 FreeSans 224 0 0 0 S2BEG[0]
port 160 nsew signal output
flabel metal2 s 18510 0 18566 56 0 FreeSans 224 0 0 0 S2BEG[1]
port 161 nsew signal output
flabel metal2 s 18786 0 18842 56 0 FreeSans 224 0 0 0 S2BEG[2]
port 162 nsew signal output
flabel metal2 s 19062 0 19118 56 0 FreeSans 224 0 0 0 S2BEG[3]
port 163 nsew signal output
flabel metal2 s 19338 0 19394 56 0 FreeSans 224 0 0 0 S2BEG[4]
port 164 nsew signal output
flabel metal2 s 19614 0 19670 56 0 FreeSans 224 0 0 0 S2BEG[5]
port 165 nsew signal output
flabel metal2 s 19890 0 19946 56 0 FreeSans 224 0 0 0 S2BEG[6]
port 166 nsew signal output
flabel metal2 s 20166 0 20222 56 0 FreeSans 224 0 0 0 S2BEG[7]
port 167 nsew signal output
flabel metal2 s 20442 0 20498 56 0 FreeSans 224 0 0 0 S2BEGb[0]
port 168 nsew signal output
flabel metal2 s 20718 0 20774 56 0 FreeSans 224 0 0 0 S2BEGb[1]
port 169 nsew signal output
flabel metal2 s 20994 0 21050 56 0 FreeSans 224 0 0 0 S2BEGb[2]
port 170 nsew signal output
flabel metal2 s 21270 0 21326 56 0 FreeSans 224 0 0 0 S2BEGb[3]
port 171 nsew signal output
flabel metal2 s 21546 0 21602 56 0 FreeSans 224 0 0 0 S2BEGb[4]
port 172 nsew signal output
flabel metal2 s 21822 0 21878 56 0 FreeSans 224 0 0 0 S2BEGb[5]
port 173 nsew signal output
flabel metal2 s 22098 0 22154 56 0 FreeSans 224 0 0 0 S2BEGb[6]
port 174 nsew signal output
flabel metal2 s 22374 0 22430 56 0 FreeSans 224 0 0 0 S2BEGb[7]
port 175 nsew signal output
flabel metal2 s 22650 0 22706 56 0 FreeSans 224 0 0 0 S4BEG[0]
port 176 nsew signal output
flabel metal2 s 25410 0 25466 56 0 FreeSans 224 0 0 0 S4BEG[10]
port 177 nsew signal output
flabel metal2 s 25686 0 25742 56 0 FreeSans 224 0 0 0 S4BEG[11]
port 178 nsew signal output
flabel metal2 s 25962 0 26018 56 0 FreeSans 224 0 0 0 S4BEG[12]
port 179 nsew signal output
flabel metal2 s 26238 0 26294 56 0 FreeSans 224 0 0 0 S4BEG[13]
port 180 nsew signal output
flabel metal2 s 26514 0 26570 56 0 FreeSans 224 0 0 0 S4BEG[14]
port 181 nsew signal output
flabel metal2 s 26790 0 26846 56 0 FreeSans 224 0 0 0 S4BEG[15]
port 182 nsew signal output
flabel metal2 s 22926 0 22982 56 0 FreeSans 224 0 0 0 S4BEG[1]
port 183 nsew signal output
flabel metal2 s 23202 0 23258 56 0 FreeSans 224 0 0 0 S4BEG[2]
port 184 nsew signal output
flabel metal2 s 23478 0 23534 56 0 FreeSans 224 0 0 0 S4BEG[3]
port 185 nsew signal output
flabel metal2 s 23754 0 23810 56 0 FreeSans 224 0 0 0 S4BEG[4]
port 186 nsew signal output
flabel metal2 s 24030 0 24086 56 0 FreeSans 224 0 0 0 S4BEG[5]
port 187 nsew signal output
flabel metal2 s 24306 0 24362 56 0 FreeSans 224 0 0 0 S4BEG[6]
port 188 nsew signal output
flabel metal2 s 24582 0 24638 56 0 FreeSans 224 0 0 0 S4BEG[7]
port 189 nsew signal output
flabel metal2 s 24858 0 24914 56 0 FreeSans 224 0 0 0 S4BEG[8]
port 190 nsew signal output
flabel metal2 s 25134 0 25190 56 0 FreeSans 224 0 0 0 S4BEG[9]
port 191 nsew signal output
flabel metal2 s 27066 0 27122 56 0 FreeSans 224 0 0 0 SS4BEG[0]
port 192 nsew signal output
flabel metal2 s 29826 0 29882 56 0 FreeSans 224 0 0 0 SS4BEG[10]
port 193 nsew signal output
flabel metal2 s 30102 0 30158 56 0 FreeSans 224 0 0 0 SS4BEG[11]
port 194 nsew signal output
flabel metal2 s 30378 0 30434 56 0 FreeSans 224 0 0 0 SS4BEG[12]
port 195 nsew signal output
flabel metal2 s 30654 0 30710 56 0 FreeSans 224 0 0 0 SS4BEG[13]
port 196 nsew signal output
flabel metal2 s 30930 0 30986 56 0 FreeSans 224 0 0 0 SS4BEG[14]
port 197 nsew signal output
flabel metal2 s 31206 0 31262 56 0 FreeSans 224 0 0 0 SS4BEG[15]
port 198 nsew signal output
flabel metal2 s 27342 0 27398 56 0 FreeSans 224 0 0 0 SS4BEG[1]
port 199 nsew signal output
flabel metal2 s 27618 0 27674 56 0 FreeSans 224 0 0 0 SS4BEG[2]
port 200 nsew signal output
flabel metal2 s 27894 0 27950 56 0 FreeSans 224 0 0 0 SS4BEG[3]
port 201 nsew signal output
flabel metal2 s 28170 0 28226 56 0 FreeSans 224 0 0 0 SS4BEG[4]
port 202 nsew signal output
flabel metal2 s 28446 0 28502 56 0 FreeSans 224 0 0 0 SS4BEG[5]
port 203 nsew signal output
flabel metal2 s 28722 0 28778 56 0 FreeSans 224 0 0 0 SS4BEG[6]
port 204 nsew signal output
flabel metal2 s 28998 0 29054 56 0 FreeSans 224 0 0 0 SS4BEG[7]
port 205 nsew signal output
flabel metal2 s 29274 0 29330 56 0 FreeSans 224 0 0 0 SS4BEG[8]
port 206 nsew signal output
flabel metal2 s 29550 0 29606 56 0 FreeSans 224 0 0 0 SS4BEG[9]
port 207 nsew signal output
flabel metal2 s 31482 0 31538 56 0 FreeSans 224 0 0 0 UserCLK
port 208 nsew signal input
flabel metal2 s 1490 11096 1546 11152 0 FreeSans 224 0 0 0 UserCLKo
port 209 nsew signal output
flabel metal4 s 3004 0 3324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 3004 11092 3324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 0 9324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 0 9324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 11092 9324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 0 15324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 0 15324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 11092 15324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 0 21324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 0 21324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 11092 21324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 0 27324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 0 27324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 11092 27324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 0 33324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 0 33324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 11092 33324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 1944 0 2264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 1944 11092 2264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 0 8264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 11092 8264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 0 14264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 0 14264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 11092 14264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 0 20264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 0 20264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 11092 20264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 0 26264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 0 26264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 11092 26264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 0 32264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 0 32264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 11092 32264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 0 38264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 0 38264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 11092 38264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
rlabel metal1 19964 8704 19964 8704 0 VGND
rlabel via1 19964 8160 19964 8160 0 VPWR
rlabel metal3 10372 1156 10372 1156 0 FrameData[0]
rlabel metal3 942 3876 942 3876 0 FrameData[10]
rlabel metal2 23322 4573 23322 4573 0 FrameData[11]
rlabel metal3 1425 4420 1425 4420 0 FrameData[12]
rlabel metal2 21390 4641 21390 4641 0 FrameData[13]
rlabel metal3 942 4964 942 4964 0 FrameData[14]
rlabel metal1 18630 4794 18630 4794 0 FrameData[15]
rlabel metal1 18814 5202 18814 5202 0 FrameData[16]
rlabel metal1 21436 5746 21436 5746 0 FrameData[17]
rlabel metal3 942 6052 942 6052 0 FrameData[18]
rlabel metal2 18722 6103 18722 6103 0 FrameData[19]
rlabel metal3 2874 1428 2874 1428 0 FrameData[1]
rlabel metal2 16698 6579 16698 6579 0 FrameData[20]
rlabel via2 15778 6851 15778 6851 0 FrameData[21]
rlabel metal3 712 7140 712 7140 0 FrameData[22]
rlabel via2 15318 7395 15318 7395 0 FrameData[23]
rlabel metal3 1425 7684 1425 7684 0 FrameData[24]
rlabel metal2 18262 7667 18262 7667 0 FrameData[25]
rlabel metal3 942 8228 942 8228 0 FrameData[26]
rlabel metal2 17066 8007 17066 8007 0 FrameData[27]
rlabel metal1 15686 7514 15686 7514 0 FrameData[28]
rlabel metal1 15778 7412 15778 7412 0 FrameData[29]
rlabel metal3 4852 1700 4852 1700 0 FrameData[2]
rlabel metal1 15456 7310 15456 7310 0 FrameData[30]
rlabel metal2 19826 8483 19826 8483 0 FrameData[31]
rlabel metal3 2920 1972 2920 1972 0 FrameData[3]
rlabel metal3 1471 2244 1471 2244 0 FrameData[4]
rlabel metal3 344 2516 344 2516 0 FrameData[5]
rlabel metal3 942 2788 942 2788 0 FrameData[6]
rlabel metal2 23046 3213 23046 3213 0 FrameData[7]
rlabel metal3 14628 3536 14628 3536 0 FrameData[8]
rlabel metal2 20746 4063 20746 4063 0 FrameData[9]
rlabel metal3 38756 1156 38756 1156 0 FrameData_O[0]
rlabel metal3 39492 3876 39492 3876 0 FrameData_O[10]
rlabel metal3 39124 4148 39124 4148 0 FrameData_O[11]
rlabel metal3 38940 4420 38940 4420 0 FrameData_O[12]
rlabel metal3 39124 4692 39124 4692 0 FrameData_O[13]
rlabel metal3 39492 4964 39492 4964 0 FrameData_O[14]
rlabel metal3 39124 5236 39124 5236 0 FrameData_O[15]
rlabel metal3 38940 5508 38940 5508 0 FrameData_O[16]
rlabel metal3 39124 5780 39124 5780 0 FrameData_O[17]
rlabel metal3 39492 6052 39492 6052 0 FrameData_O[18]
rlabel metal3 39124 6324 39124 6324 0 FrameData_O[19]
rlabel metal3 38526 1428 38526 1428 0 FrameData_O[1]
rlabel metal3 38940 6596 38940 6596 0 FrameData_O[20]
rlabel metal3 39124 6868 39124 6868 0 FrameData_O[21]
rlabel metal3 39124 7140 39124 7140 0 FrameData_O[22]
rlabel metal3 38940 7412 38940 7412 0 FrameData_O[23]
rlabel metal3 39124 7684 39124 7684 0 FrameData_O[24]
rlabel metal3 39400 7956 39400 7956 0 FrameData_O[25]
rlabel metal3 39308 8228 39308 8228 0 FrameData_O[26]
rlabel metal2 37674 8279 37674 8279 0 FrameData_O[27]
rlabel metal1 38272 7514 38272 7514 0 FrameData_O[28]
rlabel metal2 37306 8551 37306 8551 0 FrameData_O[29]
rlabel metal3 38848 1700 38848 1700 0 FrameData_O[2]
rlabel metal2 36938 8687 36938 8687 0 FrameData_O[30]
rlabel metal2 36386 9095 36386 9095 0 FrameData_O[31]
rlabel metal3 38250 1972 38250 1972 0 FrameData_O[3]
rlabel metal3 38940 2244 38940 2244 0 FrameData_O[4]
rlabel metal3 39124 2516 39124 2516 0 FrameData_O[5]
rlabel metal3 39492 2788 39492 2788 0 FrameData_O[6]
rlabel metal3 39124 3060 39124 3060 0 FrameData_O[7]
rlabel metal3 38940 3332 38940 3332 0 FrameData_O[8]
rlabel metal3 39124 3604 39124 3604 0 FrameData_O[9]
rlabel metal2 31786 3115 31786 3115 0 FrameStrobe[0]
rlabel metal2 34546 2928 34546 2928 0 FrameStrobe[10]
rlabel metal2 34822 684 34822 684 0 FrameStrobe[11]
rlabel metal2 35098 888 35098 888 0 FrameStrobe[12]
rlabel metal2 35374 2418 35374 2418 0 FrameStrobe[13]
rlabel metal2 35650 2350 35650 2350 0 FrameStrobe[14]
rlabel metal2 35926 1401 35926 1401 0 FrameStrobe[15]
rlabel metal1 35328 5746 35328 5746 0 FrameStrobe[16]
rlabel metal1 36110 5678 36110 5678 0 FrameStrobe[17]
rlabel metal1 36846 5678 36846 5678 0 FrameStrobe[18]
rlabel metal2 37030 2860 37030 2860 0 FrameStrobe[19]
rlabel metal2 32062 55 32062 55 0 FrameStrobe[1]
rlabel metal2 32338 208 32338 208 0 FrameStrobe[2]
rlabel metal1 20332 7242 20332 7242 0 FrameStrobe[3]
rlabel metal2 32890 1279 32890 1279 0 FrameStrobe[4]
rlabel metal2 33166 55 33166 55 0 FrameStrobe[5]
rlabel metal2 33442 55 33442 55 0 FrameStrobe[6]
rlabel metal2 33718 650 33718 650 0 FrameStrobe[7]
rlabel metal2 33994 3710 33994 3710 0 FrameStrobe[8]
rlabel metal2 34270 1401 34270 1401 0 FrameStrobe[9]
rlabel metal1 3680 8602 3680 8602 0 FrameStrobe_O[0]
rlabel metal1 21850 8602 21850 8602 0 FrameStrobe_O[10]
rlabel metal1 23690 8602 23690 8602 0 FrameStrobe_O[11]
rlabel metal1 25530 8602 25530 8602 0 FrameStrobe_O[12]
rlabel metal1 27416 8602 27416 8602 0 FrameStrobe_O[13]
rlabel metal1 29394 8602 29394 8602 0 FrameStrobe_O[14]
rlabel metal1 31050 8602 31050 8602 0 FrameStrobe_O[15]
rlabel metal1 32890 8602 32890 8602 0 FrameStrobe_O[16]
rlabel metal1 34730 8602 34730 8602 0 FrameStrobe_O[17]
rlabel metal1 36570 8602 36570 8602 0 FrameStrobe_O[18]
rlabel metal1 38364 8602 38364 8602 0 FrameStrobe_O[19]
rlabel metal1 5290 8602 5290 8602 0 FrameStrobe_O[1]
rlabel metal1 7130 8602 7130 8602 0 FrameStrobe_O[2]
rlabel metal1 8970 8602 8970 8602 0 FrameStrobe_O[3]
rlabel metal1 10810 8602 10810 8602 0 FrameStrobe_O[4]
rlabel metal1 12650 8602 12650 8602 0 FrameStrobe_O[5]
rlabel metal1 14490 8602 14490 8602 0 FrameStrobe_O[6]
rlabel metal1 16514 8602 16514 8602 0 FrameStrobe_O[7]
rlabel metal1 18170 8602 18170 8602 0 FrameStrobe_O[8]
rlabel metal1 20010 8602 20010 8602 0 FrameStrobe_O[9]
rlabel metal1 4094 4726 4094 4726 0 N1END[0]
rlabel metal2 3082 55 3082 55 0 N1END[1]
rlabel metal2 3358 871 3358 871 0 N1END[2]
rlabel metal1 3266 4114 3266 4114 0 N1END[3]
rlabel metal1 8326 6154 8326 6154 0 N2END[0]
rlabel metal1 8372 5814 8372 5814 0 N2END[1]
rlabel metal1 8096 6290 8096 6290 0 N2END[2]
rlabel metal1 7820 6426 7820 6426 0 N2END[3]
rlabel metal1 7728 6086 7728 6086 0 N2END[4]
rlabel metal1 7820 6698 7820 6698 0 N2END[5]
rlabel metal1 7728 6766 7728 6766 0 N2END[6]
rlabel metal2 8050 55 8050 55 0 N2END[7]
rlabel metal3 6118 5644 6118 5644 0 N2MID[0]
rlabel metal1 6900 5746 6900 5746 0 N2MID[1]
rlabel metal3 6440 4420 6440 4420 0 N2MID[2]
rlabel metal1 6026 5610 6026 5610 0 N2MID[3]
rlabel metal1 5520 5678 5520 5678 0 N2MID[4]
rlabel metal1 5014 5202 5014 5202 0 N2MID[5]
rlabel metal1 4876 5066 4876 5066 0 N2MID[6]
rlabel metal1 5152 5134 5152 5134 0 N2MID[7]
rlabel metal2 16974 3298 16974 3298 0 N4END[0]
rlabel metal1 12926 5712 12926 5712 0 N4END[10]
rlabel metal2 11362 1401 11362 1401 0 N4END[11]
rlabel metal2 11638 1347 11638 1347 0 N4END[12]
rlabel metal2 11914 1279 11914 1279 0 N4END[13]
rlabel metal1 14030 5168 14030 5168 0 N4END[14]
rlabel metal1 13524 5270 13524 5270 0 N4END[15]
rlabel metal1 17066 3060 17066 3060 0 N4END[1]
rlabel metal2 8878 55 8878 55 0 N4END[2]
rlabel metal2 9154 55 9154 55 0 N4END[3]
rlabel metal2 9430 2078 9430 2078 0 N4END[4]
rlabel metal2 9706 2316 9706 2316 0 N4END[5]
rlabel metal2 9982 1007 9982 1007 0 N4END[6]
rlabel metal1 14306 5134 14306 5134 0 N4END[7]
rlabel metal2 10534 2622 10534 2622 0 N4END[8]
rlabel metal2 10810 1500 10810 1500 0 N4END[9]
rlabel metal2 12742 191 12742 191 0 NN4END[0]
rlabel metal2 15502 1024 15502 1024 0 NN4END[10]
rlabel metal3 17319 3332 17319 3332 0 NN4END[11]
rlabel metal2 16054 276 16054 276 0 NN4END[12]
rlabel metal2 16330 939 16330 939 0 NN4END[13]
rlabel metal2 16606 174 16606 174 0 NN4END[14]
rlabel metal2 16882 871 16882 871 0 NN4END[15]
rlabel metal2 13018 140 13018 140 0 NN4END[1]
rlabel metal2 13294 327 13294 327 0 NN4END[2]
rlabel metal2 13570 259 13570 259 0 NN4END[3]
rlabel metal2 13846 106 13846 106 0 NN4END[4]
rlabel metal2 14122 55 14122 55 0 NN4END[5]
rlabel metal2 14398 55 14398 55 0 NN4END[6]
rlabel via2 14674 55 14674 55 0 NN4END[7]
rlabel metal2 14950 123 14950 123 0 NN4END[8]
rlabel metal2 15226 55 15226 55 0 NN4END[9]
rlabel metal2 17158 1160 17158 1160 0 S1BEG[0]
rlabel metal1 17572 2822 17572 2822 0 S1BEG[1]
rlabel metal2 17710 1160 17710 1160 0 S1BEG[2]
rlabel metal2 17986 1160 17986 1160 0 S1BEG[3]
rlabel metal2 18262 1160 18262 1160 0 S2BEG[0]
rlabel metal1 18676 2822 18676 2822 0 S2BEG[1]
rlabel metal2 18814 1160 18814 1160 0 S2BEG[2]
rlabel metal2 19090 1160 19090 1160 0 S2BEG[3]
rlabel metal1 19504 2822 19504 2822 0 S2BEG[4]
rlabel metal2 19642 1160 19642 1160 0 S2BEG[5]
rlabel metal2 19918 1160 19918 1160 0 S2BEG[6]
rlabel metal2 20194 1160 20194 1160 0 S2BEG[7]
rlabel metal2 20470 1160 20470 1160 0 S2BEGb[0]
rlabel metal2 20746 1160 20746 1160 0 S2BEGb[1]
rlabel metal2 21022 599 21022 599 0 S2BEGb[2]
rlabel metal2 21298 599 21298 599 0 S2BEGb[3]
rlabel metal2 21574 1296 21574 1296 0 S2BEGb[4]
rlabel metal2 21850 1330 21850 1330 0 S2BEGb[5]
rlabel metal2 22126 1194 22126 1194 0 S2BEGb[6]
rlabel metal2 22402 718 22402 718 0 S2BEGb[7]
rlabel metal1 22816 2822 22816 2822 0 S4BEG[0]
rlabel metal2 25438 1194 25438 1194 0 S4BEG[10]
rlabel metal1 25852 2822 25852 2822 0 S4BEG[11]
rlabel metal2 25990 735 25990 735 0 S4BEG[12]
rlabel metal2 26266 1296 26266 1296 0 S4BEG[13]
rlabel metal2 26542 1160 26542 1160 0 S4BEG[14]
rlabel metal2 26818 1330 26818 1330 0 S4BEG[15]
rlabel metal2 22954 1160 22954 1160 0 S4BEG[1]
rlabel metal1 23368 2822 23368 2822 0 S4BEG[2]
rlabel metal2 23506 1330 23506 1330 0 S4BEG[3]
rlabel metal1 23920 2822 23920 2822 0 S4BEG[4]
rlabel metal2 24058 1296 24058 1296 0 S4BEG[5]
rlabel metal2 24334 1194 24334 1194 0 S4BEG[6]
rlabel metal2 24610 1330 24610 1330 0 S4BEG[7]
rlabel metal1 25024 2822 25024 2822 0 S4BEG[8]
rlabel metal2 25162 1296 25162 1296 0 S4BEG[9]
rlabel metal2 27094 55 27094 55 0 SS4BEG[0]
rlabel metal2 29854 1330 29854 1330 0 SS4BEG[10]
rlabel metal2 30130 1296 30130 1296 0 SS4BEG[11]
rlabel metal1 30544 2822 30544 2822 0 SS4BEG[12]
rlabel metal2 30682 1296 30682 1296 0 SS4BEG[13]
rlabel metal1 31096 2822 31096 2822 0 SS4BEG[14]
rlabel metal2 31234 599 31234 599 0 SS4BEG[15]
rlabel metal2 27370 1296 27370 1296 0 SS4BEG[1]
rlabel metal2 27646 1194 27646 1194 0 SS4BEG[2]
rlabel metal2 27922 599 27922 599 0 SS4BEG[3]
rlabel metal1 28290 2822 28290 2822 0 SS4BEG[4]
rlabel metal1 28612 2822 28612 2822 0 SS4BEG[5]
rlabel metal2 28750 1296 28750 1296 0 SS4BEG[6]
rlabel metal2 29026 1160 29026 1160 0 SS4BEG[7]
rlabel metal1 29394 2822 29394 2822 0 SS4BEG[8]
rlabel metal2 29578 1058 29578 1058 0 SS4BEG[9]
rlabel metal2 31510 735 31510 735 0 UserCLK
rlabel metal1 1564 8602 1564 8602 0 UserCLKo
rlabel metal1 37490 2448 37490 2448 0 net1
rlabel metal2 17802 5814 17802 5814 0 net10
rlabel metal1 28934 3060 28934 3060 0 net100
rlabel metal1 30636 2278 30636 2278 0 net101
rlabel metal1 30268 3910 30268 3910 0 net102
rlabel metal1 30038 3026 30038 3026 0 net103
rlabel metal1 30176 2482 30176 2482 0 net104
rlabel metal1 1794 8500 1794 8500 0 net105
rlabel metal2 19090 6120 19090 6120 0 net11
rlabel metal2 36846 2142 36846 2142 0 net12
rlabel metal1 18584 6426 18584 6426 0 net13
rlabel metal2 16146 6749 16146 6749 0 net14
rlabel metal2 20194 6528 20194 6528 0 net15
rlabel metal2 15686 7548 15686 7548 0 net16
rlabel metal2 18814 7514 18814 7514 0 net17
rlabel metal1 18446 7310 18446 7310 0 net18
rlabel metal2 19734 7786 19734 7786 0 net19
rlabel metal1 37858 4182 37858 4182 0 net2
rlabel metal1 21666 7344 21666 7344 0 net20
rlabel metal1 21758 7412 21758 7412 0 net21
rlabel metal2 15962 7072 15962 7072 0 net22
rlabel metal2 37490 3536 37490 3536 0 net23
rlabel metal2 16882 7718 16882 7718 0 net24
rlabel metal2 36202 8840 36202 8840 0 net25
rlabel metal2 32246 2244 32246 2244 0 net26
rlabel metal1 37858 2482 37858 2482 0 net27
rlabel metal2 38226 2210 38226 2210 0 net28
rlabel metal1 37858 3094 37858 3094 0 net29
rlabel metal2 38226 4420 38226 4420 0 net3
rlabel metal2 37950 3230 37950 3230 0 net30
rlabel metal1 34799 3502 34799 3502 0 net31
rlabel via2 22034 3995 22034 3995 0 net32
rlabel metal2 21850 7599 21850 7599 0 net33
rlabel metal1 25162 5882 25162 5882 0 net34
rlabel metal2 28842 6426 28842 6426 0 net35
rlabel metal1 26956 3978 26956 3978 0 net36
rlabel metal1 28612 4794 28612 4794 0 net37
rlabel metal2 30774 6630 30774 6630 0 net38
rlabel metal2 31326 6902 31326 6902 0 net39
rlabel metal1 31050 4556 31050 4556 0 net4
rlabel metal2 34270 7174 34270 7174 0 net40
rlabel metal1 35282 5882 35282 5882 0 net41
rlabel metal1 36800 5882 36800 5882 0 net42
rlabel metal1 37398 5882 37398 5882 0 net43
rlabel metal1 17894 7174 17894 7174 0 net44
rlabel metal1 21160 7174 21160 7174 0 net45
rlabel metal1 17158 7242 17158 7242 0 net46
rlabel metal2 17250 8772 17250 8772 0 net47
rlabel metal2 12926 8772 12926 8772 0 net48
rlabel metal2 14766 8806 14766 8806 0 net49
rlabel metal1 38226 4556 38226 4556 0 net5
rlabel metal2 16974 8670 16974 8670 0 net50
rlabel metal2 18446 8636 18446 8636 0 net51
rlabel metal1 20286 8500 20286 8500 0 net52
rlabel metal1 16192 2414 16192 2414 0 net53
rlabel metal1 17526 2958 17526 2958 0 net54
rlabel metal2 17342 3876 17342 3876 0 net55
rlabel metal1 17710 2380 17710 2380 0 net56
rlabel metal2 18078 1870 18078 1870 0 net57
rlabel metal3 14812 3332 14812 3332 0 net58
rlabel metal1 18446 2482 18446 2482 0 net59
rlabel metal1 37858 5236 37858 5236 0 net6
rlabel metal2 18814 4318 18814 4318 0 net60
rlabel metal2 12742 5848 12742 5848 0 net61
rlabel metal2 8602 6358 8602 6358 0 net62
rlabel metal2 19642 2482 19642 2482 0 net63
rlabel metal1 19734 2448 19734 2448 0 net64
rlabel metal1 20424 2414 20424 2414 0 net65
rlabel metal2 20562 1989 20562 1989 0 net66
rlabel metal2 20838 2142 20838 2142 0 net67
rlabel metal1 18354 2414 18354 2414 0 net68
rlabel metal2 9982 6137 9982 6137 0 net69
rlabel metal2 19642 4930 19642 4930 0 net7
rlabel metal2 22310 2176 22310 2176 0 net70
rlabel metal3 12489 2380 12489 2380 0 net71
rlabel metal1 23184 2414 23184 2414 0 net72
rlabel metal2 17618 3944 17618 3944 0 net73
rlabel metal2 25990 2074 25990 2074 0 net74
rlabel metal1 21942 3944 21942 3944 0 net75
rlabel metal1 16606 3604 16606 3604 0 net76
rlabel metal1 26220 2482 26220 2482 0 net77
rlabel metal2 17986 3230 17986 3230 0 net78
rlabel metal1 19044 3638 19044 3638 0 net79
rlabel metal1 20286 5338 20286 5338 0 net8
rlabel metal2 14490 2213 14490 2213 0 net80
rlabel metal2 21574 4250 21574 4250 0 net81
rlabel metal2 13386 3672 13386 3672 0 net82
rlabel metal2 23874 3536 23874 3536 0 net83
rlabel metal2 13110 3808 13110 3808 0 net84
rlabel metal1 20838 2550 20838 2550 0 net85
rlabel metal2 13846 4828 13846 4828 0 net86
rlabel metal1 14490 5100 14490 5100 0 net87
rlabel metal1 19274 4488 19274 4488 0 net88
rlabel metal2 27462 3468 27462 3468 0 net89
rlabel metal1 38226 5644 38226 5644 0 net9
rlabel metal1 30636 2414 30636 2414 0 net90
rlabel metal1 29900 3706 29900 3706 0 net91
rlabel metal1 30544 3026 30544 3026 0 net92
rlabel metal1 29670 5134 29670 5134 0 net93
rlabel metal1 31050 2992 31050 2992 0 net94
rlabel metal2 32154 2108 32154 2108 0 net95
rlabel metal1 28014 2414 28014 2414 0 net96
rlabel metal1 28796 2414 28796 2414 0 net97
rlabel metal1 29026 2414 29026 2414 0 net98
rlabel metal1 28704 3026 28704 3026 0 net99
<< properties >>
string FIXED_BBOX 0 0 39928 11152
<< end >>
