module RAM_IO (Config_accessC_bit0,
    Config_accessC_bit1,
    Config_accessC_bit2,
    Config_accessC_bit3,
    FAB2RAM_A0_O0,
    FAB2RAM_A0_O1,
    FAB2RAM_A0_O2,
    FAB2RAM_A0_O3,
    FAB2RAM_A1_O0,
    FAB2RAM_A1_O1,
    FAB2RAM_A1_O2,
    FAB2RAM_A1_O3,
    FAB2RAM_C_O0,
    FAB2RAM_C_O1,
    FAB2RAM_C_O2,
    FAB2RAM_C_O3,
    FAB2RAM_D0_O0,
    FAB2RAM_D0_O1,
    FAB2RAM_D0_O2,
    FAB2RAM_D0_O3,
    FAB2RAM_D1_O0,
    FAB2RAM_D1_O1,
    FAB2RAM_D1_O2,
    FAB2RAM_D1_O3,
    FAB2RAM_D2_O0,
    FAB2RAM_D2_O1,
    FAB2RAM_D2_O2,
    FAB2RAM_D2_O3,
    FAB2RAM_D3_O0,
    FAB2RAM_D3_O1,
    FAB2RAM_D3_O2,
    FAB2RAM_D3_O3,
    RAM2FAB_D0_I0,
    RAM2FAB_D0_I1,
    RAM2FAB_D0_I2,
    RAM2FAB_D0_I3,
    RAM2FAB_D1_I0,
    RAM2FAB_D1_I1,
    RAM2FAB_D1_I2,
    RAM2FAB_D1_I3,
    RAM2FAB_D2_I0,
    RAM2FAB_D2_I1,
    RAM2FAB_D2_I2,
    RAM2FAB_D2_I3,
    RAM2FAB_D3_I0,
    RAM2FAB_D3_I1,
    RAM2FAB_D3_I2,
    RAM2FAB_D3_I3,
    UserCLK,
    UserCLKo,
    VGND,
    VPWR,
    E1END,
    E2END,
    E2MID,
    E6END,
    EE4END,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N1END,
    N2BEG,
    N2BEGb,
    N2END,
    N2MID,
    N4BEG,
    N4END,
    S1BEG,
    S1END,
    S2BEG,
    S2BEGb,
    S2END,
    S2MID,
    S4BEG,
    S4END,
    W1BEG,
    W2BEG,
    W2BEGb,
    W6BEG,
    WW4BEG);
 output Config_accessC_bit0;
 output Config_accessC_bit1;
 output Config_accessC_bit2;
 output Config_accessC_bit3;
 output FAB2RAM_A0_O0;
 output FAB2RAM_A0_O1;
 output FAB2RAM_A0_O2;
 output FAB2RAM_A0_O3;
 output FAB2RAM_A1_O0;
 output FAB2RAM_A1_O1;
 output FAB2RAM_A1_O2;
 output FAB2RAM_A1_O3;
 output FAB2RAM_C_O0;
 output FAB2RAM_C_O1;
 output FAB2RAM_C_O2;
 output FAB2RAM_C_O3;
 output FAB2RAM_D0_O0;
 output FAB2RAM_D0_O1;
 output FAB2RAM_D0_O2;
 output FAB2RAM_D0_O3;
 output FAB2RAM_D1_O0;
 output FAB2RAM_D1_O1;
 output FAB2RAM_D1_O2;
 output FAB2RAM_D1_O3;
 output FAB2RAM_D2_O0;
 output FAB2RAM_D2_O1;
 output FAB2RAM_D2_O2;
 output FAB2RAM_D2_O3;
 output FAB2RAM_D3_O0;
 output FAB2RAM_D3_O1;
 output FAB2RAM_D3_O2;
 output FAB2RAM_D3_O3;
 input RAM2FAB_D0_I0;
 input RAM2FAB_D0_I1;
 input RAM2FAB_D0_I2;
 input RAM2FAB_D0_I3;
 input RAM2FAB_D1_I0;
 input RAM2FAB_D1_I1;
 input RAM2FAB_D1_I2;
 input RAM2FAB_D1_I3;
 input RAM2FAB_D2_I0;
 input RAM2FAB_D2_I1;
 input RAM2FAB_D2_I2;
 input RAM2FAB_D2_I3;
 input RAM2FAB_D3_I0;
 input RAM2FAB_D3_I1;
 input RAM2FAB_D3_I2;
 input RAM2FAB_D3_I3;
 input UserCLK;
 output UserCLKo;
 input VGND;
 input VPWR;
 input [3:0] E1END;
 input [7:0] E2END;
 input [7:0] E2MID;
 input [11:0] E6END;
 input [15:0] EE4END;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 input [3:0] N1END;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 input [7:0] N2END;
 input [7:0] N2MID;
 output [15:0] N4BEG;
 input [15:0] N4END;
 output [3:0] S1BEG;
 input [3:0] S1END;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 input [7:0] S2END;
 input [7:0] S2MID;
 output [15:0] S4BEG;
 input [15:0] S4END;
 output [3:0] W1BEG;
 output [7:0] W2BEG;
 output [7:0] W2BEGb;
 output [11:0] W6BEG;
 output [15:0] WW4BEG;

 wire \Inst_Config_accessConfig_access.ConfigBits[0] ;
 wire \Inst_Config_accessConfig_access.ConfigBits[1] ;
 wire \Inst_Config_accessConfig_access.ConfigBits[2] ;
 wire \Inst_Config_accessConfig_access.ConfigBits[3] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits[0] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits[1] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits[2] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits[3] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I[0] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I[1] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I[2] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I[3] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q[0] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q[1] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q[2] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q[3] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._0_ ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._1_ ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._0_ ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._1_ ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._0_ ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._1_ ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._0_ ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._1_ ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits[0] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits[1] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits[2] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits[3] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I[0] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I[1] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I[2] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I[3] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q[0] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q[1] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q[2] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q[3] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._0_ ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._1_ ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._0_ ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._1_ ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._0_ ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._1_ ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._0_ ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._1_ ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits[0] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits[1] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits[2] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits[3] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.I[0] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.I[1] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.I[2] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.I[3] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q[0] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q[1] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q[2] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q[3] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._0_ ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._1_ ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._0_ ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._1_ ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._0_ ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._1_ ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._0_ ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._1_ ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits[0] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits[1] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits[2] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits[3] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I[0] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I[1] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I[2] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I[3] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q[0] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q[1] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q[2] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q[3] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._0_ ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._1_ ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._0_ ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._1_ ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._0_ ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._1_ ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._0_ ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._1_ ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits[0] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits[1] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits[2] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits[3] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I[0] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I[1] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I[2] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I[3] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q[0] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q[1] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q[2] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q[3] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._0_ ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._1_ ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._0_ ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._1_ ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._0_ ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._1_ ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._0_ ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._1_ ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits[0] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits[1] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits[2] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits[3] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I[0] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I[1] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I[2] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I[3] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q[0] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q[1] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q[2] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q[3] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._0_ ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._1_ ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._0_ ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._1_ ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._0_ ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._1_ ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._0_ ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._1_ ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits[0] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits[1] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits[2] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits[3] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I[0] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I[1] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I[2] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I[3] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q[0] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q[1] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q[2] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q[3] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._0_ ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._1_ ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._0_ ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._1_ ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._0_ ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._1_ ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._0_ ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._1_ ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits[0] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits[1] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits[2] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits[3] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[0] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[1] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[2] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[3] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q[0] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q[1] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q[2] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q[3] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._0_ ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._1_ ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._0_ ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._1_ ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._0_ ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._1_ ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._0_ ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._1_ ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits[0] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits[1] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits[2] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits[3] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[0] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[1] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[2] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[3] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q[0] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q[1] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q[2] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q[3] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._0_ ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._1_ ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._0_ ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._1_ ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._0_ ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._1_ ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._0_ ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._1_ ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits[0] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits[1] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits[2] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits[3] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[0] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[1] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[2] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[3] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q[0] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q[1] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q[2] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q[3] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._0_ ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._1_ ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._0_ ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._1_ ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._0_ ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._1_ ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._0_ ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._1_ ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits[0] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits[1] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits[2] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits[3] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[0] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[1] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[2] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[3] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q[0] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q[1] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q[2] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q[3] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._0_ ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._1_ ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._0_ ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._1_ ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._0_ ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._1_ ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._0_ ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._1_ ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[100] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[101] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[102] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[103] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[104] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[105] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[106] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[107] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[108] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[109] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[110] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[111] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[112] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[113] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[114] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[115] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[116] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[117] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[118] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[119] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[120] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[121] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[122] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[123] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[124] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[125] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[126] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[127] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[128] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[129] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[130] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[131] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[132] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[133] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[134] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[135] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[136] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[137] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[138] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[139] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[140] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[141] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[142] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[143] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[144] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[145] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[146] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[147] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[148] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[149] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[150] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[151] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[152] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[153] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[154] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[155] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[156] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[157] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[158] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[159] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[160] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[161] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[162] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[163] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[164] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[165] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[166] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[167] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[168] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[169] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[170] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[171] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[172] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[173] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[174] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[175] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[176] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[177] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[178] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[179] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[180] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[181] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[182] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[183] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[184] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[185] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[186] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[187] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[188] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[189] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[190] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[191] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[192] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[193] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[194] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[195] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[196] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[197] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[198] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[199] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[200] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[201] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[202] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[203] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[204] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[205] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[206] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[207] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[208] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[209] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[210] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[211] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[212] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[213] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[214] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[215] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[216] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[217] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[218] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[219] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[220] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[221] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[222] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[223] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[224] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[225] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[226] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[227] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[228] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[229] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[230] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[231] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[232] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[233] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[234] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[235] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[236] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[237] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[238] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[239] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[240] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[241] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[242] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[243] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[244] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[245] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[246] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[247] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[248] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[249] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[250] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[251] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[252] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[253] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[254] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[255] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[256] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[257] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[258] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[259] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[260] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[261] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[262] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[263] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[264] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[265] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[266] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[267] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[268] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[269] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[270] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[271] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[272] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[273] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[274] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[275] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[276] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[277] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[278] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[279] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[280] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[281] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[282] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[283] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[284] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[285] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[286] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[287] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[288] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[289] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[290] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[291] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[292] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[293] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[294] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[295] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[296] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[297] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[298] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[299] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[300] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[301] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[302] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[303] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[304] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[305] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[306] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[307] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[308] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[309] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[310] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[311] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[312] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[313] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[314] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[315] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[316] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[317] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[318] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[319] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[320] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[321] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[322] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[323] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[324] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[325] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[326] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[327] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[48] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[49] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[50] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[51] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[52] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[53] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[54] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[55] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[56] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[57] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[58] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[59] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[60] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[61] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[62] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[63] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[64] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[65] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[66] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[67] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[68] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[69] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[70] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[71] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[72] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[73] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[74] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[75] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[76] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[77] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[78] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[79] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[80] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[81] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[82] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[83] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[84] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[85] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[86] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[87] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[88] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[89] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[90] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[91] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[92] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[93] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[94] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[95] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[96] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[97] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[98] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits[99] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[0] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[100] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[101] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[102] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[103] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[104] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[105] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[106] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[107] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[108] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[109] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[10] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[110] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[111] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[112] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[113] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[114] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[115] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[116] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[117] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[118] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[119] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[11] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[120] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[121] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[122] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[123] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[124] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[125] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[126] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[127] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[128] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[129] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[12] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[130] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[131] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[132] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[133] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[134] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[135] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[136] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[137] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[138] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[139] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[13] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[140] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[141] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[142] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[143] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[144] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[145] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[146] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[147] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[148] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[149] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[14] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[150] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[151] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[152] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[153] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[154] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[155] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[156] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[157] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[158] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[159] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[15] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[160] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[161] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[162] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[163] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[164] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[165] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[166] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[167] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[168] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[169] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[16] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[170] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[171] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[172] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[173] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[174] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[175] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[176] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[177] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[178] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[179] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[17] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[180] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[181] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[182] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[183] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[184] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[185] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[186] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[187] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[188] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[189] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[18] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[190] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[191] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[192] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[193] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[194] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[195] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[196] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[197] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[198] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[199] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[19] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[1] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[200] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[201] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[202] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[203] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[204] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[205] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[206] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[207] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[208] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[209] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[20] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[210] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[211] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[212] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[213] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[214] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[215] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[216] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[217] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[218] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[219] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[21] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[220] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[221] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[222] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[223] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[224] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[225] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[226] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[227] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[228] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[229] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[22] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[230] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[231] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[232] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[233] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[234] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[235] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[236] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[237] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[238] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[239] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[23] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[240] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[241] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[242] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[243] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[244] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[245] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[246] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[247] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[248] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[249] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[24] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[250] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[251] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[252] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[253] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[254] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[255] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[256] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[257] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[258] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[259] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[25] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[260] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[261] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[262] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[263] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[264] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[265] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[266] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[267] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[268] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[269] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[26] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[270] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[271] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[272] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[273] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[274] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[275] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[276] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[277] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[278] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[279] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[27] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[280] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[281] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[282] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[283] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[284] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[285] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[286] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[287] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[288] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[289] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[28] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[290] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[291] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[292] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[293] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[294] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[295] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[296] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[297] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[298] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[299] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[29] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[2] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[300] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[301] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[302] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[303] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[304] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[305] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[306] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[307] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[308] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[309] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[30] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[310] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[311] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[312] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[313] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[314] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[315] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[316] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[317] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[318] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[319] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[31] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[320] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[321] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[322] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[323] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[324] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[325] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[326] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[327] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[32] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[33] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[34] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[35] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[36] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[37] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[38] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[39] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[3] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[40] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[41] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[42] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[43] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[44] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[45] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[46] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[47] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[48] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[49] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[4] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[50] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[51] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[52] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[53] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[54] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[55] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[56] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[57] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[58] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[59] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[5] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[60] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[61] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[62] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[63] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[64] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[65] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[66] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[67] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[68] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[69] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[6] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[70] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[71] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[72] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[73] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[74] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[75] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[76] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[77] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[78] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[79] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[7] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[80] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[81] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[82] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[83] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[84] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[85] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[86] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[87] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[88] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[89] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[8] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[90] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[91] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[92] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[93] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[94] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[95] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[96] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[97] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[98] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[99] ;
 wire \Inst_RAM_IO_ConfigMem.ConfigBits_N[9] ;
 wire \Inst_RAM_IO_switch_matrix.J_NS1_BEG0 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS1_BEG1 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS1_BEG2 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS1_BEG3 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS2_BEG0 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS2_BEG1 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS2_BEG2 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS2_BEG3 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS2_BEG4 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS2_BEG5 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS2_BEG6 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS2_BEG7 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS4_BEG0 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS4_BEG1 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS4_BEG10 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS4_BEG11 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS4_BEG12 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS4_BEG13 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS4_BEG14 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS4_BEG15 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS4_BEG2 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS4_BEG3 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS4_BEG4 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS4_BEG5 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS4_BEG6 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS4_BEG7 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS4_BEG8 ;
 wire \Inst_RAM_IO_switch_matrix.J_NS4_BEG9 ;
 wire \Inst_RAM_IO_switch_matrix.N1BEG0 ;
 wire \Inst_RAM_IO_switch_matrix.N1BEG1 ;
 wire \Inst_RAM_IO_switch_matrix.N1BEG2 ;
 wire \Inst_RAM_IO_switch_matrix.N1BEG3 ;
 wire \Inst_RAM_IO_switch_matrix.N2BEG0 ;
 wire \Inst_RAM_IO_switch_matrix.N2BEG1 ;
 wire \Inst_RAM_IO_switch_matrix.N2BEG2 ;
 wire \Inst_RAM_IO_switch_matrix.N2BEG3 ;
 wire \Inst_RAM_IO_switch_matrix.N2BEG4 ;
 wire \Inst_RAM_IO_switch_matrix.N2BEG5 ;
 wire \Inst_RAM_IO_switch_matrix.N2BEG6 ;
 wire \Inst_RAM_IO_switch_matrix.N2BEG7 ;
 wire \Inst_RAM_IO_switch_matrix.N2BEGb0 ;
 wire \Inst_RAM_IO_switch_matrix.N2BEGb1 ;
 wire \Inst_RAM_IO_switch_matrix.N2BEGb2 ;
 wire \Inst_RAM_IO_switch_matrix.N2BEGb3 ;
 wire \Inst_RAM_IO_switch_matrix.N2BEGb4 ;
 wire \Inst_RAM_IO_switch_matrix.N2BEGb5 ;
 wire \Inst_RAM_IO_switch_matrix.N2BEGb6 ;
 wire \Inst_RAM_IO_switch_matrix.N2BEGb7 ;
 wire \Inst_RAM_IO_switch_matrix.N4BEG0 ;
 wire \Inst_RAM_IO_switch_matrix.N4BEG1 ;
 wire \Inst_RAM_IO_switch_matrix.N4BEG2 ;
 wire \Inst_RAM_IO_switch_matrix.N4BEG3 ;
 wire \Inst_RAM_IO_switch_matrix.S1BEG0 ;
 wire \Inst_RAM_IO_switch_matrix.S1BEG1 ;
 wire \Inst_RAM_IO_switch_matrix.S1BEG2 ;
 wire \Inst_RAM_IO_switch_matrix.S1BEG3 ;
 wire \Inst_RAM_IO_switch_matrix.S2BEG0 ;
 wire \Inst_RAM_IO_switch_matrix.S2BEG1 ;
 wire \Inst_RAM_IO_switch_matrix.S2BEG2 ;
 wire \Inst_RAM_IO_switch_matrix.S2BEG3 ;
 wire \Inst_RAM_IO_switch_matrix.S2BEG4 ;
 wire \Inst_RAM_IO_switch_matrix.S2BEG5 ;
 wire \Inst_RAM_IO_switch_matrix.S2BEG6 ;
 wire \Inst_RAM_IO_switch_matrix.S2BEG7 ;
 wire \Inst_RAM_IO_switch_matrix.S2BEGb0 ;
 wire \Inst_RAM_IO_switch_matrix.S2BEGb1 ;
 wire \Inst_RAM_IO_switch_matrix.S2BEGb2 ;
 wire \Inst_RAM_IO_switch_matrix.S2BEGb3 ;
 wire \Inst_RAM_IO_switch_matrix.S2BEGb4 ;
 wire \Inst_RAM_IO_switch_matrix.S2BEGb5 ;
 wire \Inst_RAM_IO_switch_matrix.S2BEGb6 ;
 wire \Inst_RAM_IO_switch_matrix.S2BEGb7 ;
 wire \Inst_RAM_IO_switch_matrix.S4BEG0 ;
 wire \Inst_RAM_IO_switch_matrix.S4BEG1 ;
 wire \Inst_RAM_IO_switch_matrix.S4BEG2 ;
 wire \Inst_RAM_IO_switch_matrix.S4BEG3 ;
 wire \Inst_RAM_IO_switch_matrix.W1BEG0 ;
 wire \Inst_RAM_IO_switch_matrix.W1BEG1 ;
 wire \Inst_RAM_IO_switch_matrix.W1BEG2 ;
 wire \Inst_RAM_IO_switch_matrix.W1BEG3 ;
 wire \Inst_RAM_IO_switch_matrix.W2BEG0 ;
 wire \Inst_RAM_IO_switch_matrix.W2BEG1 ;
 wire \Inst_RAM_IO_switch_matrix.W2BEG2 ;
 wire \Inst_RAM_IO_switch_matrix.W2BEG3 ;
 wire \Inst_RAM_IO_switch_matrix.W2BEG4 ;
 wire \Inst_RAM_IO_switch_matrix.W2BEG5 ;
 wire \Inst_RAM_IO_switch_matrix.W2BEG6 ;
 wire \Inst_RAM_IO_switch_matrix.W2BEG7 ;
 wire \Inst_RAM_IO_switch_matrix.W2BEGb0 ;
 wire \Inst_RAM_IO_switch_matrix.W2BEGb1 ;
 wire \Inst_RAM_IO_switch_matrix.W2BEGb2 ;
 wire \Inst_RAM_IO_switch_matrix.W2BEGb3 ;
 wire \Inst_RAM_IO_switch_matrix.W2BEGb4 ;
 wire \Inst_RAM_IO_switch_matrix.W2BEGb5 ;
 wire \Inst_RAM_IO_switch_matrix.W2BEGb6 ;
 wire \Inst_RAM_IO_switch_matrix.W2BEGb7 ;
 wire \Inst_RAM_IO_switch_matrix.W6BEG0 ;
 wire \Inst_RAM_IO_switch_matrix.W6BEG1 ;
 wire \Inst_RAM_IO_switch_matrix.W6BEG10 ;
 wire \Inst_RAM_IO_switch_matrix.W6BEG11 ;
 wire \Inst_RAM_IO_switch_matrix.W6BEG2 ;
 wire \Inst_RAM_IO_switch_matrix.W6BEG3 ;
 wire \Inst_RAM_IO_switch_matrix.W6BEG4 ;
 wire \Inst_RAM_IO_switch_matrix.W6BEG5 ;
 wire \Inst_RAM_IO_switch_matrix.W6BEG6 ;
 wire \Inst_RAM_IO_switch_matrix.W6BEG7 ;
 wire \Inst_RAM_IO_switch_matrix.W6BEG8 ;
 wire \Inst_RAM_IO_switch_matrix.W6BEG9 ;
 wire \Inst_RAM_IO_switch_matrix.WW4BEG0 ;
 wire \Inst_RAM_IO_switch_matrix.WW4BEG1 ;
 wire \Inst_RAM_IO_switch_matrix.WW4BEG10 ;
 wire \Inst_RAM_IO_switch_matrix.WW4BEG11 ;
 wire \Inst_RAM_IO_switch_matrix.WW4BEG12 ;
 wire \Inst_RAM_IO_switch_matrix.WW4BEG13 ;
 wire \Inst_RAM_IO_switch_matrix.WW4BEG14 ;
 wire \Inst_RAM_IO_switch_matrix.WW4BEG15 ;
 wire \Inst_RAM_IO_switch_matrix.WW4BEG2 ;
 wire \Inst_RAM_IO_switch_matrix.WW4BEG3 ;
 wire \Inst_RAM_IO_switch_matrix.WW4BEG4 ;
 wire \Inst_RAM_IO_switch_matrix.WW4BEG5 ;
 wire \Inst_RAM_IO_switch_matrix.WW4BEG6 ;
 wire \Inst_RAM_IO_switch_matrix.WW4BEG7 ;
 wire \Inst_RAM_IO_switch_matrix.WW4BEG8 ;
 wire \Inst_RAM_IO_switch_matrix.WW4BEG9 ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.A0 ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.A1 ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.AIN[0] ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.AIN[1] ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._0_ ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._1_ ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.A0 ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.A1 ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.AIN[0] ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.AIN[1] ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._0_ ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._1_ ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.A0 ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.A1 ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.AIN[0] ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.AIN[1] ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._0_ ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._1_ ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.A0 ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.A1 ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.AIN[0] ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.AIN[1] ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._0_ ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._1_ ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.A0 ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.A1 ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.AIN[0] ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.AIN[1] ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._0_ ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._1_ ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.A0 ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.A1 ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.AIN[0] ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.AIN[1] ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._0_ ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._1_ ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.A0 ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.A1 ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.AIN[0] ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.AIN[1] ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._0_ ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._1_ ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.A0 ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.A1 ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.AIN[0] ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.AIN[1] ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._0_ ;
 wire \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._1_ ;
 wire \N4BEG_outbuf_0.A ;
 wire \N4BEG_outbuf_0.X ;
 wire \N4BEG_outbuf_1.A ;
 wire \N4BEG_outbuf_1.X ;
 wire \N4BEG_outbuf_10.A ;
 wire \N4BEG_outbuf_10.X ;
 wire \N4BEG_outbuf_11.A ;
 wire \N4BEG_outbuf_11.X ;
 wire \N4BEG_outbuf_2.A ;
 wire \N4BEG_outbuf_2.X ;
 wire \N4BEG_outbuf_3.A ;
 wire \N4BEG_outbuf_3.X ;
 wire \N4BEG_outbuf_4.A ;
 wire \N4BEG_outbuf_4.X ;
 wire \N4BEG_outbuf_5.A ;
 wire \N4BEG_outbuf_5.X ;
 wire \N4BEG_outbuf_6.A ;
 wire \N4BEG_outbuf_6.X ;
 wire \N4BEG_outbuf_7.A ;
 wire \N4BEG_outbuf_7.X ;
 wire \N4BEG_outbuf_8.A ;
 wire \N4BEG_outbuf_8.X ;
 wire \N4BEG_outbuf_9.A ;
 wire \N4BEG_outbuf_9.X ;
 wire \S4BEG_outbuf_0.A ;
 wire \S4BEG_outbuf_0.X ;
 wire \S4BEG_outbuf_1.A ;
 wire \S4BEG_outbuf_1.X ;
 wire \S4BEG_outbuf_10.A ;
 wire \S4BEG_outbuf_10.X ;
 wire \S4BEG_outbuf_11.A ;
 wire \S4BEG_outbuf_11.X ;
 wire \S4BEG_outbuf_2.A ;
 wire \S4BEG_outbuf_2.X ;
 wire \S4BEG_outbuf_3.A ;
 wire \S4BEG_outbuf_3.X ;
 wire \S4BEG_outbuf_4.A ;
 wire \S4BEG_outbuf_4.X ;
 wire \S4BEG_outbuf_5.A ;
 wire \S4BEG_outbuf_5.X ;
 wire \S4BEG_outbuf_6.A ;
 wire \S4BEG_outbuf_6.X ;
 wire \S4BEG_outbuf_7.A ;
 wire \S4BEG_outbuf_7.X ;
 wire \S4BEG_outbuf_8.A ;
 wire \S4BEG_outbuf_8.X ;
 wire \S4BEG_outbuf_9.A ;
 wire \S4BEG_outbuf_9.X ;
 wire \data_inbuf_0.X ;
 wire \data_inbuf_1.X ;
 wire \data_inbuf_10.X ;
 wire \data_inbuf_11.X ;
 wire \data_inbuf_12.X ;
 wire \data_inbuf_13.X ;
 wire \data_inbuf_14.X ;
 wire \data_inbuf_15.X ;
 wire \data_inbuf_16.X ;
 wire \data_inbuf_17.X ;
 wire \data_inbuf_18.X ;
 wire \data_inbuf_19.X ;
 wire \data_inbuf_2.X ;
 wire \data_inbuf_20.X ;
 wire \data_inbuf_21.X ;
 wire \data_inbuf_22.X ;
 wire \data_inbuf_23.X ;
 wire \data_inbuf_24.X ;
 wire \data_inbuf_25.X ;
 wire \data_inbuf_26.X ;
 wire \data_inbuf_27.X ;
 wire \data_inbuf_28.X ;
 wire \data_inbuf_29.X ;
 wire \data_inbuf_3.X ;
 wire \data_inbuf_30.X ;
 wire \data_inbuf_31.X ;
 wire \data_inbuf_4.X ;
 wire \data_inbuf_5.X ;
 wire \data_inbuf_6.X ;
 wire \data_inbuf_7.X ;
 wire \data_inbuf_8.X ;
 wire \data_inbuf_9.X ;
 wire \data_outbuf_0.X ;
 wire \data_outbuf_1.X ;
 wire \data_outbuf_10.X ;
 wire \data_outbuf_11.X ;
 wire \data_outbuf_12.X ;
 wire \data_outbuf_13.X ;
 wire \data_outbuf_14.X ;
 wire \data_outbuf_15.X ;
 wire \data_outbuf_16.X ;
 wire \data_outbuf_17.X ;
 wire \data_outbuf_18.X ;
 wire \data_outbuf_19.X ;
 wire \data_outbuf_2.X ;
 wire \data_outbuf_20.X ;
 wire \data_outbuf_21.X ;
 wire \data_outbuf_22.X ;
 wire \data_outbuf_23.X ;
 wire \data_outbuf_24.X ;
 wire \data_outbuf_25.X ;
 wire \data_outbuf_26.X ;
 wire \data_outbuf_27.X ;
 wire \data_outbuf_28.X ;
 wire \data_outbuf_29.X ;
 wire \data_outbuf_3.X ;
 wire \data_outbuf_30.X ;
 wire \data_outbuf_31.X ;
 wire \data_outbuf_4.X ;
 wire \data_outbuf_5.X ;
 wire \data_outbuf_6.X ;
 wire \data_outbuf_7.X ;
 wire \data_outbuf_8.X ;
 wire \data_outbuf_9.X ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \strobe_inbuf_0.X ;
 wire \strobe_inbuf_1.X ;
 wire \strobe_inbuf_10.X ;
 wire \strobe_inbuf_11.X ;
 wire \strobe_inbuf_12.X ;
 wire \strobe_inbuf_13.X ;
 wire \strobe_inbuf_14.X ;
 wire \strobe_inbuf_15.X ;
 wire \strobe_inbuf_16.X ;
 wire \strobe_inbuf_17.X ;
 wire \strobe_inbuf_18.X ;
 wire \strobe_inbuf_19.X ;
 wire \strobe_inbuf_2.X ;
 wire \strobe_inbuf_3.X ;
 wire \strobe_inbuf_4.X ;
 wire \strobe_inbuf_5.X ;
 wire \strobe_inbuf_6.X ;
 wire \strobe_inbuf_7.X ;
 wire \strobe_inbuf_8.X ;
 wire \strobe_inbuf_9.X ;
 wire \strobe_outbuf_0.X ;
 wire \strobe_outbuf_1.X ;
 wire \strobe_outbuf_10.X ;
 wire \strobe_outbuf_11.X ;
 wire \strobe_outbuf_12.X ;
 wire \strobe_outbuf_13.X ;
 wire \strobe_outbuf_14.X ;
 wire \strobe_outbuf_15.X ;
 wire \strobe_outbuf_16.X ;
 wire \strobe_outbuf_17.X ;
 wire \strobe_outbuf_18.X ;
 wire \strobe_outbuf_19.X ;
 wire \strobe_outbuf_2.X ;
 wire \strobe_outbuf_3.X ;
 wire \strobe_outbuf_4.X ;
 wire \strobe_outbuf_5.X ;
 wire \strobe_outbuf_6.X ;
 wire \strobe_outbuf_7.X ;
 wire \strobe_outbuf_8.X ;
 wire \strobe_outbuf_9.X ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(FrameStrobe[19]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\Inst_RAM_IO_switch_matrix.S2BEG4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\Inst_RAM_IO_switch_matrix.S2BEGb4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(RAM2FAB_D1_I1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\S4BEG_outbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\S4BEG_outbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\Inst_RAM_IO_switch_matrix.S2BEG5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\strobe_inbuf_16.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\S4BEG_outbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net349),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(\S4BEG_outbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(\S4BEG_outbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\Inst_RAM_IO_switch_matrix.S2BEGb7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\N4BEG_outbuf_3.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\N4BEG_outbuf_5.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(RAM2FAB_D0_I1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(RAM2FAB_D1_I3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\strobe_inbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_40_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_43_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_44_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_44_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_44_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_45_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_45_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_45_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_47_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_47_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_48_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_49_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_51_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_53_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_54_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_56_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_56_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_57_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_57_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_57_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_57_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_58_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_58_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_59_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_61_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_61_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_63_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_63_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_63_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_64_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_66_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_66_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_66_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_67_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_67_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_67_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_67_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_67_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_67_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_68_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_69_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_74_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_1 \Inst_Config_accessConfig_access._0_  (.A(\Inst_Config_accessConfig_access.ConfigBits[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 \Inst_Config_accessConfig_access._1_  (.A(\Inst_Config_accessConfig_access.ConfigBits[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 \Inst_Config_accessConfig_access._2_  (.A(\Inst_Config_accessConfig_access.ConfigBits[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 \Inst_Config_accessConfig_access._3_  (.A(\Inst_Config_accessConfig_access.ConfigBits[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net192));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux._0_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux._1_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux._2_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux._3_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._2_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._3_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ),
    .B(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._4_  (.A1(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits[0] ),
    .A2(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._0_ ),
    .B1(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net193));
 sky130_fd_sc_hd__buf_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._2_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._3_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ),
    .B(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._4_  (.A1(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits[1] ),
    .A2(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._0_ ),
    .B1(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net194));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._2_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._3_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ),
    .B(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._4_  (.A1(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits[2] ),
    .A2(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._0_ ),
    .B1(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net195));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._2_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._3_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ),
    .B(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._4_  (.A1(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits[3] ),
    .A2(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._0_ ),
    .B1(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net196));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux._0_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux._1_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux._2_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux._3_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._2_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._3_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ),
    .B(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._4_  (.A1(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits[0] ),
    .A2(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._0_ ),
    .B1(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net197));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._2_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._3_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ),
    .B(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._4_  (.A1(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits[1] ),
    .A2(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._0_ ),
    .B1(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net198));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._2_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._3_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ),
    .B(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._4_  (.A1(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits[2] ),
    .A2(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._0_ ),
    .B1(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net199));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._2_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._3_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ),
    .B(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._4_  (.A1(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits[3] ),
    .A2(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._0_ ),
    .B1(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net200));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux._0_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux._1_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux._2_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux._3_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._2_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._3_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ),
    .B(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._4_  (.A1(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits[0] ),
    .A2(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._0_ ),
    .B1(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net201));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._2_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._3_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ),
    .B(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._4_  (.A1(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits[1] ),
    .A2(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._0_ ),
    .B1(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net202));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._2_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._3_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ),
    .B(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._4_  (.A1(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits[2] ),
    .A2(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._0_ ),
    .B1(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net203));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._2_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._3_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ),
    .B(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._4_  (.A1(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits[3] ),
    .A2(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._0_ ),
    .B1(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net204));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux._0_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux._1_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux._2_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux._3_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._2_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._3_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ),
    .B(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._4_  (.A1(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits[0] ),
    .A2(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._0_ ),
    .B1(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net205));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._2_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._3_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ),
    .B(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._4_  (.A1(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits[1] ),
    .A2(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._0_ ),
    .B1(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net206));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._2_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._3_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ),
    .B(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._4_  (.A1(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits[2] ),
    .A2(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._0_ ),
    .B1(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net207));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._2_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._3_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ),
    .B(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._4_  (.A1(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits[3] ),
    .A2(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._0_ ),
    .B1(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net208));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux._0_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux._1_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux._2_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux._3_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._2_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._3_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ),
    .B(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._4_  (.A1(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits[0] ),
    .A2(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._0_ ),
    .B1(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net209));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._2_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._3_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ),
    .B(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._4_  (.A1(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits[1] ),
    .A2(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._0_ ),
    .B1(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net210));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._2_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._3_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ),
    .B(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._4_  (.A1(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits[2] ),
    .A2(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._0_ ),
    .B1(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net211));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._2_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._3_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ),
    .B(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._4_  (.A1(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits[3] ),
    .A2(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._0_ ),
    .B1(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net212));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux._0_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux._1_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux._2_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux._3_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._2_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._3_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ),
    .B(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._4_  (.A1(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits[0] ),
    .A2(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._0_ ),
    .B1(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net213));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._2_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._3_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ),
    .B(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._4_  (.A1(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits[1] ),
    .A2(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._0_ ),
    .B1(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net214));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._2_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._3_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ),
    .B(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._4_  (.A1(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits[2] ),
    .A2(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._0_ ),
    .B1(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net215));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._2_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._3_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ),
    .B(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._4_  (.A1(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits[3] ),
    .A2(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._0_ ),
    .B1(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net216));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux._0_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux._1_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux._2_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux._3_  (.CLK(UserCLK),
    .D(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._2_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._3_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ),
    .B(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._4_  (.A1(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits[0] ),
    .A2(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._0_ ),
    .B1(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net217));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._2_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._3_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ),
    .B(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._4_  (.A1(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits[1] ),
    .A2(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._0_ ),
    .B1(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net218));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._2_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._3_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ),
    .B(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._4_  (.A1(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits[2] ),
    .A2(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._0_ ),
    .B1(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net219));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._2_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._3_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ),
    .B(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._4_  (.A1(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits[3] ),
    .A2(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._0_ ),
    .B1(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net220));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux._0_  (.CLK(UserCLK),
    .D(net137),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux._1_  (.CLK(UserCLK),
    .D(net138),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux._2_  (.CLK(UserCLK),
    .D(net139),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux._3_  (.CLK(UserCLK),
    .D(net140),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._2_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._3_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ),
    .B(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._4_  (.A1(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits[0] ),
    .A2(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._0_ ),
    .B1(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_  (.A(net137),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._2_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._3_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ),
    .B(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._4_  (.A1(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits[1] ),
    .A2(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._0_ ),
    .B1(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[1] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_  (.A(net138),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._2_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._3_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ),
    .B(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._4_  (.A1(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits[2] ),
    .A2(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._0_ ),
    .B1(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[2] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_  (.A(net139),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._2_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._3_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ),
    .B(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._4_  (.A1(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits[3] ),
    .A2(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._0_ ),
    .B1(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[3] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_  (.A(net140),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux._0_  (.CLK(UserCLK),
    .D(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux._1_  (.CLK(UserCLK),
    .D(net142),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux._2_  (.CLK(UserCLK),
    .D(net143),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux._3_  (.CLK(UserCLK),
    .D(net144),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._2_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._3_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ),
    .B(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._4_  (.A1(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits[0] ),
    .A2(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._0_ ),
    .B1(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_  (.A(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._2_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._3_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ),
    .B(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._4_  (.A1(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits[1] ),
    .A2(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._0_ ),
    .B1(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[1] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_  (.A(net142),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._2_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._3_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ),
    .B(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._4_  (.A1(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits[2] ),
    .A2(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._0_ ),
    .B1(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[2] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_  (.A(net143),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._2_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._3_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ),
    .B(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._4_  (.A1(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits[3] ),
    .A2(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._0_ ),
    .B1(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[3] ));
 sky130_fd_sc_hd__buf_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_  (.A(net144),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux._0_  (.CLK(UserCLK),
    .D(net145),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux._1_  (.CLK(UserCLK),
    .D(net146),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux._2_  (.CLK(UserCLK),
    .D(net147),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux._3_  (.CLK(UserCLK),
    .D(net148),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._2_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._3_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ),
    .B(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._4_  (.A1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits[0] ),
    .A2(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._0_ ),
    .B1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_  (.A(net145),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._2_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._3_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ),
    .B(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._4_  (.A1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits[1] ),
    .A2(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._0_ ),
    .B1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[1] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_  (.A(net146),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._2_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._3_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ),
    .B(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._4_  (.A1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits[2] ),
    .A2(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._0_ ),
    .B1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[2] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_  (.A(net147),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._2_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._3_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ),
    .B(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._4_  (.A1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits[3] ),
    .A2(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._0_ ),
    .B1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[3] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_  (.A(net148),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux._0_  (.CLK(UserCLK),
    .D(net149),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux._1_  (.CLK(UserCLK),
    .D(net150),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux._2_  (.CLK(UserCLK),
    .D(net151),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux._3_  (.CLK(UserCLK),
    .D(net152),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._2_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._3_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ),
    .B(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._4_  (.A1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits[0] ),
    .A2(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._0_ ),
    .B1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_  (.A(net149),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._2_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._3_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ),
    .B(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._4_  (.A1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits[1] ),
    .A2(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._0_ ),
    .B1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[1] ));
 sky130_fd_sc_hd__buf_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_  (.A(net150),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._2_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._3_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ),
    .B(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._4_  (.A1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits[2] ),
    .A2(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._0_ ),
    .B1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[2] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_  (.A(net151),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._2_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._3_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ),
    .B(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._4_  (.A1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits[3] ),
    .A2(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._0_ ),
    .B1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[3] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_  (.A(net152),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.AIN[1] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit0  (.D(net49),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[296] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[296] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit1  (.D(net60),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[297] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[297] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit10  (.D(net50),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[306] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[306] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit11  (.D(net51),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[307] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[307] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit12  (.D(net52),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[308] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[308] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit13  (.D(net53),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[309] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[309] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit14  (.D(net54),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[310] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[310] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit15  (.D(net55),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[311] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[311] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit16  (.D(net56),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[312] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[312] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit17  (.D(net57),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[313] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[313] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit18  (.D(net58),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[314] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[314] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit19  (.D(net59),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[315] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[315] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit2  (.D(net71),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[298] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[298] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit20  (.D(net61),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[316] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[316] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit21  (.D(net62),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[317] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[317] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit22  (.D(net63),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[318] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[318] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit23  (.D(net64),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[319] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[319] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit24  (.D(net65),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[320] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[320] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit25  (.D(net66),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[321] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[321] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit26  (.D(net67),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[322] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[322] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit27  (.D(net68),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[323] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[323] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit28  (.D(net69),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[324] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[324] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit29  (.D(net70),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[325] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[325] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit3  (.D(net74),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[299] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[299] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit30  (.D(net72),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[326] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[326] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit31  (.D(net73),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[327] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[327] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit4  (.D(net75),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[300] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[300] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit5  (.D(net76),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[301] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[301] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit6  (.D(net77),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[302] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[302] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit7  (.D(net78),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[303] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[303] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit8  (.D(net79),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[304] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[304] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame0_bit9  (.D(net80),
    .GATE(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[305] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[305] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame10_bit24  (.D(net65),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits[0] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[0] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame10_bit25  (.D(net66),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits[1] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[1] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame10_bit26  (.D(net67),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits[2] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[2] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame10_bit27  (.D(net68),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits[3] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[3] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame10_bit28  (.D(net69),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits[0] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[4] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame10_bit29  (.D(net70),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits[1] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[5] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame10_bit30  (.D(net72),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits[2] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[6] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame10_bit31  (.D(net73),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits[3] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[7] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit0  (.D(net49),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[264] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[264] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit1  (.D(net60),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[265] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[265] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit10  (.D(net50),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[274] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[274] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit11  (.D(net51),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[275] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[275] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit12  (.D(net52),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[276] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[276] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit13  (.D(net53),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[277] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[277] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit14  (.D(net54),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[278] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[278] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit15  (.D(net55),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[279] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[279] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit16  (.D(net56),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[280] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[280] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit17  (.D(net57),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[281] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[281] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit18  (.D(net58),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[282] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[282] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit19  (.D(net59),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[283] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[283] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit2  (.D(net71),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[266] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[266] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit20  (.D(net61),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[284] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[284] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit21  (.D(net62),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[285] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[285] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit22  (.D(net63),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[286] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[286] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit23  (.D(net64),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[287] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[287] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit24  (.D(net65),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[288] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[288] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit25  (.D(net66),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[289] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[289] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit26  (.D(net67),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[290] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[290] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit27  (.D(net68),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[291] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[291] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit28  (.D(net69),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[292] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[292] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit29  (.D(net70),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[293] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[293] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit3  (.D(net74),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[267] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[267] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit30  (.D(net72),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[294] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[294] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit31  (.D(net73),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[295] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[295] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit4  (.D(net75),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[268] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[268] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit5  (.D(net76),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[269] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[269] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit6  (.D(net77),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[270] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[270] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit7  (.D(net78),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[271] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[271] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit8  (.D(net79),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[272] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[272] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame1_bit9  (.D(net80),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[273] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[273] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit0  (.D(net49),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[232] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[232] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit1  (.D(net60),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[233] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[233] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit10  (.D(net50),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[242] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[242] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit11  (.D(net51),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[243] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[243] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit12  (.D(net52),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[244] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[244] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit13  (.D(net53),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[245] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[245] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit14  (.D(net54),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[246] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[246] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit15  (.D(net55),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[247] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[247] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit16  (.D(net56),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[248] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[248] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit17  (.D(net57),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[249] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[249] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit18  (.D(net58),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[250] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[250] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit19  (.D(net59),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[251] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[251] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit2  (.D(net71),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[234] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[234] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit20  (.D(net61),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[252] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[252] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit21  (.D(net62),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[253] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[253] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit22  (.D(net63),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[254] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[254] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit23  (.D(net64),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[255] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[255] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit24  (.D(net65),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[256] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[256] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit25  (.D(net66),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[257] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[257] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit26  (.D(net67),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[258] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[258] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit27  (.D(net68),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[259] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[259] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit28  (.D(net69),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[260] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[260] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit29  (.D(net70),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[261] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[261] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit3  (.D(net74),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[235] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[235] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit30  (.D(net72),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[262] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[262] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit31  (.D(net73),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[263] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[263] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit4  (.D(net75),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[236] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[236] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit5  (.D(net76),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[237] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[237] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit6  (.D(net77),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[238] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[238] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit7  (.D(net78),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[239] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[239] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit8  (.D(net79),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[240] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[240] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame2_bit9  (.D(net80),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[241] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[241] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit0  (.D(net49),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[200] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[200] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit1  (.D(net60),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[201] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[201] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit10  (.D(net50),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[210] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[210] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit11  (.D(net51),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[211] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[211] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit12  (.D(net52),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[212] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[212] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit13  (.D(net53),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[213] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[213] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit14  (.D(net54),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[214] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[214] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit15  (.D(net55),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[215] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[215] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit16  (.D(net56),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[216] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[216] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit17  (.D(net57),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[217] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[217] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit18  (.D(net58),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[218] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[218] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit19  (.D(net59),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[219] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[219] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit2  (.D(net71),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[202] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[202] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit20  (.D(net61),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[220] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[220] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit21  (.D(net62),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[221] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[221] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit22  (.D(net63),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[222] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[222] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit23  (.D(net64),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[223] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[223] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit24  (.D(net65),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[224] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[224] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit25  (.D(net66),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[225] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[225] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit26  (.D(net67),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[226] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[226] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit27  (.D(net68),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[227] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[227] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit28  (.D(net69),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[228] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[228] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit29  (.D(net70),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[229] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[229] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit3  (.D(net74),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[203] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[203] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit30  (.D(net72),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[230] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[230] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit31  (.D(net73),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[231] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[231] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit4  (.D(net75),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[204] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[204] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit5  (.D(net76),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[205] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[205] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit6  (.D(net77),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[206] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[206] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit7  (.D(net78),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[207] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[207] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit8  (.D(net79),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[208] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[208] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame3_bit9  (.D(net80),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[209] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[209] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit0  (.D(net49),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[168] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[168] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit1  (.D(net60),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[169] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[169] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit10  (.D(net50),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[178] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[178] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit11  (.D(net51),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[179] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[179] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit12  (.D(net52),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[180] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[180] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit13  (.D(net53),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[181] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[181] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit14  (.D(net54),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[182] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[182] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit15  (.D(net55),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[183] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[183] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit16  (.D(net56),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[184] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[184] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit17  (.D(net57),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[185] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[185] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit18  (.D(net58),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[186] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[186] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit19  (.D(net59),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[187] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[187] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit2  (.D(net71),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[170] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[170] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit20  (.D(net61),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[188] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[188] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit21  (.D(net62),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[189] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[189] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit22  (.D(net63),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[190] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[190] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit23  (.D(net64),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[191] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[191] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit24  (.D(net65),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[192] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[192] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit25  (.D(net66),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[193] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[193] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit26  (.D(net67),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[194] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[194] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit27  (.D(net68),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[195] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[195] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit28  (.D(net69),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[196] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[196] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit29  (.D(net70),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[197] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[197] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit3  (.D(net74),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[171] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[171] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit30  (.D(net72),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[198] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[198] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit31  (.D(net73),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[199] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[199] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit4  (.D(net75),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[172] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[172] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit5  (.D(net76),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[173] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[173] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit6  (.D(net77),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[174] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[174] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit7  (.D(net78),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[175] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[175] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit8  (.D(net79),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[176] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[176] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame4_bit9  (.D(net80),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[177] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[177] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit0  (.D(net49),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[136] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[136] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit1  (.D(net60),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[137] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[137] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit10  (.D(net50),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[146] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[146] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit11  (.D(net51),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[147] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[147] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit12  (.D(net52),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[148] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[148] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit13  (.D(net53),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[149] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[149] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit14  (.D(net54),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[150] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[150] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit15  (.D(net55),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[151] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[151] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit16  (.D(net56),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[152] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[152] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit17  (.D(net57),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[153] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[153] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit18  (.D(net58),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[154] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[154] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit19  (.D(net59),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[155] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[155] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit2  (.D(net71),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[138] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[138] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit20  (.D(net61),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[156] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[156] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit21  (.D(net62),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[157] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[157] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit22  (.D(net63),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[158] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[158] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit23  (.D(net64),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[159] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[159] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit24  (.D(net65),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[160] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[160] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit25  (.D(net66),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[161] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[161] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit26  (.D(net67),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[162] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[162] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit27  (.D(net68),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[163] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[163] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit28  (.D(net69),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[164] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[164] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit29  (.D(net70),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[165] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[165] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit3  (.D(net74),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[139] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[139] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit30  (.D(net72),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[166] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[166] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit31  (.D(net73),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[167] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[167] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit4  (.D(net75),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[140] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[140] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit5  (.D(net76),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[141] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[141] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit6  (.D(net77),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[142] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[142] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit7  (.D(net78),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[143] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[143] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit8  (.D(net79),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[144] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[144] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame5_bit9  (.D(net80),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[145] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[145] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit0  (.D(net49),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[104] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[104] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit1  (.D(net60),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[105] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[105] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit10  (.D(net50),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[114] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[114] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit11  (.D(net51),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[115] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[115] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit12  (.D(net52),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[116] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[116] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit13  (.D(net53),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[117] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[117] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit14  (.D(net54),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[118] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[118] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit15  (.D(net55),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[119] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[119] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit16  (.D(net56),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[120] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[120] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit17  (.D(net57),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[121] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[121] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit18  (.D(net58),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[122] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[122] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit19  (.D(net59),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[123] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[123] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit2  (.D(net71),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[106] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[106] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit20  (.D(net61),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[124] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[124] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit21  (.D(net62),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[125] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[125] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit22  (.D(net63),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[126] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[126] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit23  (.D(net64),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[127] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[127] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit24  (.D(net65),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[128] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[128] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit25  (.D(net66),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[129] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[129] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit26  (.D(net67),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[130] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[130] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit27  (.D(net68),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[131] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[131] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit28  (.D(net69),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[132] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[132] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit29  (.D(net70),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[133] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[133] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit3  (.D(net74),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[107] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[107] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit30  (.D(net72),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[134] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[134] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit31  (.D(net73),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[135] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[135] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit4  (.D(net75),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[108] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[108] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit5  (.D(net76),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[109] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[109] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit6  (.D(net77),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[110] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[110] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit7  (.D(net78),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[111] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[111] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit8  (.D(net79),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[112] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[112] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame6_bit9  (.D(net80),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[113] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[113] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit0  (.D(net49),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[72] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[72] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit1  (.D(net60),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[73] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[73] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit10  (.D(net50),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[82] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[82] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit11  (.D(net51),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[83] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[83] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit12  (.D(net52),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[84] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[84] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit13  (.D(net53),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[85] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[85] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit14  (.D(net54),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[86] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[86] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit15  (.D(net55),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[87] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[87] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit16  (.D(net56),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[88] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[88] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit17  (.D(net57),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[89] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[89] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit18  (.D(net58),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[90] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[90] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit19  (.D(net59),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[91] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[91] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit2  (.D(net71),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[74] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[74] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit20  (.D(net61),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[92] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[92] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit21  (.D(net62),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[93] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[93] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit22  (.D(net63),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[94] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[94] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit23  (.D(net64),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[95] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[95] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit24  (.D(net65),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[96] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[96] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit25  (.D(net66),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[97] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[97] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit26  (.D(net67),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[98] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[98] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit27  (.D(net68),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[99] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[99] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit28  (.D(net69),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[100] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[100] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit29  (.D(net70),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[101] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[101] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit3  (.D(net74),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[75] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[75] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit30  (.D(net72),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[102] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[102] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit31  (.D(net73),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[103] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[103] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit4  (.D(net75),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[76] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[76] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit5  (.D(net76),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[77] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[77] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit6  (.D(net77),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[78] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[78] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit7  (.D(net78),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[79] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[79] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit8  (.D(net79),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[80] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[80] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame7_bit9  (.D(net80),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[81] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[81] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit0  (.D(net49),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits[0] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[40] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit1  (.D(net60),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits[1] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[41] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit10  (.D(net50),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[50] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[50] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit11  (.D(net51),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[51] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[51] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit12  (.D(net52),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[52] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[52] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit13  (.D(net53),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[53] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[53] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit14  (.D(net54),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[54] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[54] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit15  (.D(net55),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[55] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[55] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit16  (.D(net56),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[56] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[56] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit17  (.D(net57),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[57] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[57] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit18  (.D(net58),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[58] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[58] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit19  (.D(net59),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[59] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[59] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit2  (.D(net71),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits[2] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[42] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit20  (.D(net61),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[60] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[60] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit21  (.D(net62),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[61] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[61] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit22  (.D(net63),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[62] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[62] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit23  (.D(net64),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[63] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[63] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit24  (.D(net65),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[64] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[64] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit25  (.D(net66),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[65] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[65] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit26  (.D(net67),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[66] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[66] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit27  (.D(net68),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[67] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[67] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit28  (.D(net69),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[68] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[68] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit29  (.D(net70),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[69] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[69] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit3  (.D(net74),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits[3] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[43] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit30  (.D(net72),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[70] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[70] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit31  (.D(net73),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[71] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[71] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit4  (.D(net75),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_Config_accessConfig_access.ConfigBits[0] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[44] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit5  (.D(net76),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_Config_accessConfig_access.ConfigBits[1] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[45] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit6  (.D(net77),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_Config_accessConfig_access.ConfigBits[2] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[46] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit7  (.D(net78),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_Config_accessConfig_access.ConfigBits[3] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[47] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit8  (.D(net79),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[48] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[48] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame8_bit9  (.D(net80),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM_IO_ConfigMem.ConfigBits[49] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[49] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit0  (.D(net49),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits[0] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[8] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit1  (.D(net60),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits[1] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[9] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit10  (.D(net50),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits[2] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[18] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit11  (.D(net51),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits[3] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[19] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit12  (.D(net52),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits[0] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[20] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit13  (.D(net53),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits[1] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[21] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit14  (.D(net54),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits[2] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[22] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit15  (.D(net55),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits[3] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[23] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit16  (.D(net56),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits[0] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[24] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit17  (.D(net57),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits[1] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[25] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit18  (.D(net58),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits[2] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[26] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit19  (.D(net59),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits[3] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[27] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit2  (.D(net71),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits[2] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[10] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit20  (.D(net61),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits[0] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[28] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit21  (.D(net62),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits[1] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[29] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit22  (.D(net63),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits[2] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[30] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit23  (.D(net64),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits[3] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[31] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit24  (.D(net65),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits[0] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[32] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit25  (.D(net66),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits[1] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[33] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit26  (.D(net67),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits[2] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[34] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit27  (.D(net68),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits[3] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[35] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit28  (.D(net69),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits[0] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[36] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit29  (.D(net70),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits[1] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[37] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit3  (.D(net74),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits[3] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[11] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit30  (.D(net72),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits[2] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[38] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit31  (.D(net73),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits[3] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[39] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit4  (.D(net75),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits[0] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[12] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit5  (.D(net76),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits[1] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[13] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit6  (.D(net77),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits[2] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[14] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit7  (.D(net78),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits[3] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[15] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit8  (.D(net79),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits[0] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[16] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem.Inst_frame9_bit9  (.D(net80),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits[1] ),
    .Q_N(\Inst_RAM_IO_ConfigMem.ConfigBits_N[17] ));
 sky130_fd_sc_hd__buf_1 \Inst_RAM_IO_switch_matrix._32_  (.A(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.N2BEGb0 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix._33_  (.A(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.N2BEGb1 ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RAM_IO_switch_matrix._34_  (.A(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.N2BEGb2 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix._35_  (.A(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.N2BEGb3 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix._36_  (.A(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.N2BEGb4 ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RAM_IO_switch_matrix._37_  (.A(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.N2BEGb5 ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RAM_IO_switch_matrix._38_  (.A(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.N2BEGb6 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix._39_  (.A(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.N2BEGb7 ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RAM_IO_switch_matrix._40_  (.A(net165),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.S2BEGb0 ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RAM_IO_switch_matrix._41_  (.A(net166),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.S2BEGb1 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix._42_  (.A(net167),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.S2BEGb2 ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RAM_IO_switch_matrix._43_  (.A(net168),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.S2BEGb3 ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RAM_IO_switch_matrix._44_  (.A(net169),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.S2BEGb4 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix._45_  (.A(net170),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.S2BEGb5 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix._46_  (.A(net171),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.S2BEGb6 ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RAM_IO_switch_matrix._47_  (.A(net172),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.S2BEGb7 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I0  (.A0(net13),
    .A1(net5),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG0 ),
    .A3(net395),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[248] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[249] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I[0] ));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I0_395  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net395));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I1  (.A0(net14),
    .A1(net6),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG1 ),
    .A3(net396),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[250] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[251] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I[1] ));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I1_396  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net396));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I2  (.A0(net15),
    .A1(net7),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG2 ),
    .A3(net397),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[252] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[253] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I[2] ));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I2_397  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net397));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I3  (.A0(net16),
    .A1(net8),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG3 ),
    .A3(net398),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[254] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[255] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I[3] ));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I3_398  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net398));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I0  (.A0(net17),
    .A1(net9),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG4 ),
    .A3(net399),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[256] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[257] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I[0] ));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I0_399  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net399));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I1  (.A0(net18),
    .A1(net10),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG5 ),
    .A3(net400),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[258] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[259] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I[1] ));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I1_400  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net400));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I2  (.A0(net19),
    .A1(net11),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG6 ),
    .A3(net401),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[260] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[261] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I[2] ));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I2_401  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net401));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I3  (.A0(net20),
    .A1(net12),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG7 ),
    .A3(net402),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[262] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[263] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I[3] ));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I3_402  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net402));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I0  (.A0(net1),
    .A1(net21),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS1_BEG0 ),
    .A3(net403),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[264] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[265] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.I[0] ));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I0_403  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net403));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I1  (.A0(net2),
    .A1(net24),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS1_BEG1 ),
    .A3(net404),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[266] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[267] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.I[1] ));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I1_404  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net404));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I2  (.A0(net3),
    .A1(net25),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS1_BEG2 ),
    .A3(net405),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[268] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[269] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.I[2] ));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I2_405  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net405));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I3  (.A0(net4),
    .A1(net26),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS1_BEG3 ),
    .A3(net409),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[270] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[271] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_C_OutPass4_frame_config_mux.I[3] ));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I3_409  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net409));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I0  (.A0(net33),
    .A1(net47),
    .A2(net21),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG0 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[216] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[217] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I1  (.A0(net40),
    .A1(net48),
    .A2(net24),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG1 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[218] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[219] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I2  (.A0(net41),
    .A1(net34),
    .A2(net25),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG2 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[220] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[221] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I3  (.A0(net42),
    .A1(net35),
    .A2(net26),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG3 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[222] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[223] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I0  (.A0(net43),
    .A1(net36),
    .A2(net27),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG4 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[224] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[225] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I1  (.A0(net44),
    .A1(net37),
    .A2(net28),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG5 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[226] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[227] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I2  (.A0(net45),
    .A1(net38),
    .A2(net29),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG6 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[228] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[229] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I3  (.A0(net46),
    .A1(net39),
    .A2(net30),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG7 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[230] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[231] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I[3] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I0  (.A0(net33),
    .A1(net47),
    .A2(net31),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG8 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[232] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[233] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I1  (.A0(net40),
    .A1(net48),
    .A2(net32),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG9 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[234] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[235] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I2  (.A0(net41),
    .A1(net34),
    .A2(net22),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG10 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[236] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[237] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I3  (.A0(net42),
    .A1(net35),
    .A2(net23),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG11 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[238] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[239] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I0  (.A0(net1),
    .A1(net43),
    .A2(net36),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG12 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[240] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[241] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I1  (.A0(net2),
    .A1(net44),
    .A2(net37),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG13 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[242] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[243] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I2  (.A0(net3),
    .A1(net45),
    .A2(net38),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG14 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[244] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[245] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I3  (.A0(net4),
    .A1(net46),
    .A2(net39),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG15 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[246] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[247] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I[3] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG0  (.A0(net101),
    .A1(net21),
    .A2(net153),
    .A3(net406),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[320] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[321] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS1_BEG0 ));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG0_406  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net406));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG1  (.A0(net102),
    .A1(net24),
    .A2(net154),
    .A3(net407),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[322] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[323] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS1_BEG1 ));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG1_407  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net407));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG2  (.A0(net103),
    .A1(net25),
    .A2(net155),
    .A3(net408),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[324] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[325] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS1_BEG2 ));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG2_408  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net408));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG3  (.A0(net104),
    .A1(net26),
    .A2(net156),
    .A3(net394),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[326] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[327] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS1_BEG3 ));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG3_394  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net394));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG0  (.A0(net113),
    .A1(net105),
    .A2(net165),
    .A3(net157),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[304] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[305] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS2_BEG0 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG1  (.A0(net114),
    .A1(net106),
    .A2(net166),
    .A3(net158),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[306] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[307] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS2_BEG1 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG2  (.A0(net115),
    .A1(net107),
    .A2(net167),
    .A3(net159),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[308] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[309] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS2_BEG2 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG3  (.A0(net116),
    .A1(net108),
    .A2(net168),
    .A3(net160),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[310] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[311] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS2_BEG3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG4  (.A0(net117),
    .A1(net109),
    .A2(net169),
    .A3(net161),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[312] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[313] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS2_BEG4 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG5  (.A0(net118),
    .A1(net110),
    .A2(net170),
    .A3(net162),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[314] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[315] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS2_BEG5 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG6  (.A0(net119),
    .A1(net111),
    .A2(net171),
    .A3(net163),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[316] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[317] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS2_BEG6 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG7  (.A0(net120),
    .A1(net112),
    .A2(net172),
    .A3(net164),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[318] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[319] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS2_BEG7 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG0  (.A0(net101),
    .A1(net121),
    .A2(net153),
    .A3(net173),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[272] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[273] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS4_BEG0 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG1  (.A0(net102),
    .A1(net128),
    .A2(net154),
    .A3(net180),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[274] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[275] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS4_BEG1 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG10  (.A0(net103),
    .A1(net129),
    .A2(net155),
    .A3(net181),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[292] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[293] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS4_BEG10 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG11  (.A0(net104),
    .A1(net130),
    .A2(net156),
    .A3(net182),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[294] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[295] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS4_BEG11 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG12  (.A0(net101),
    .A1(net121),
    .A2(net153),
    .A3(net173),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[296] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[297] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS4_BEG12 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG13  (.A0(net102),
    .A1(net128),
    .A2(net154),
    .A3(net180),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[298] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[299] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS4_BEG13 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG14  (.A0(net103),
    .A1(net129),
    .A2(net155),
    .A3(net181),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[300] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[301] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS4_BEG14 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG15  (.A0(net104),
    .A1(net130),
    .A2(net156),
    .A3(net182),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[302] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[303] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS4_BEG15 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG2  (.A0(net103),
    .A1(net129),
    .A2(net155),
    .A3(net181),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[276] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[277] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS4_BEG2 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG3  (.A0(net104),
    .A1(net130),
    .A2(net156),
    .A3(net182),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[278] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[279] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS4_BEG3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG4  (.A0(net101),
    .A1(net121),
    .A2(net153),
    .A3(net173),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[280] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[281] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS4_BEG4 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG5  (.A0(net102),
    .A1(net128),
    .A2(net154),
    .A3(net180),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[282] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[283] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS4_BEG5 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG6  (.A0(net103),
    .A1(net129),
    .A2(net155),
    .A3(net181),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[284] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[285] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS4_BEG6 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG7  (.A0(net104),
    .A1(net130),
    .A2(net156),
    .A3(net182),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[286] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[287] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS4_BEG7 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG8  (.A0(net101),
    .A1(net121),
    .A2(net153),
    .A3(net173),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[288] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[289] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS4_BEG8 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG9  (.A0(net102),
    .A1(net128),
    .A2(net154),
    .A3(net180),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[290] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[291] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.J_NS4_BEG9 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG0  (.A0(net1),
    .A1(net27),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG12 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS1_BEG0 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[48] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.N1BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG1  (.A0(net2),
    .A1(net28),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG13 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS1_BEG1 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[50] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.N1BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG2  (.A0(net3),
    .A1(net29),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG14 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS1_BEG2 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[52] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.N1BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG3  (.A0(net4),
    .A1(net30),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG15 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS1_BEG3 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[54] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.N1BEG3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG0  (.A0(net20),
    .A1(net12),
    .A2(net30),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG0 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[56] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.N2BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG1  (.A0(net19),
    .A1(net11),
    .A2(net29),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG1 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[58] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.N2BEG1 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG2  (.A0(net18),
    .A1(net10),
    .A2(net28),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG2 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[60] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.N2BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG3  (.A0(net17),
    .A1(net9),
    .A2(net27),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG3 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[62] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.N2BEG3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG4  (.A0(net16),
    .A1(net8),
    .A2(net26),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG4 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[64] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.N2BEG4 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG5  (.A0(net15),
    .A1(net7),
    .A2(net25),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG5 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[66] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.N2BEG5 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG6  (.A0(net14),
    .A1(net6),
    .A2(net24),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG6 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[68] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.N2BEG6 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG7  (.A0(net13),
    .A1(net5),
    .A2(net21),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG7 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[70] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.N2BEG7 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG0  (.A0(net1),
    .A1(net31),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG12 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS1_BEG0 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[84] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.S1BEG0 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG1  (.A0(net2),
    .A1(net32),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG13 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS1_BEG1 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[86] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.S1BEG1 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG2  (.A0(net3),
    .A1(net22),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG14 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS1_BEG2 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[88] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.S1BEG2 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG3  (.A0(net4),
    .A1(net23),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG15 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS1_BEG3 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[90] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.S1BEG3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG0  (.A0(net20),
    .A1(net12),
    .A2(net31),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG0 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[92] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.S2BEG0 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG1  (.A0(net19),
    .A1(net11),
    .A2(net32),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG1 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[94] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.S2BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG2  (.A0(net18),
    .A1(net10),
    .A2(net22),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG2 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[96] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.S2BEG2 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG3  (.A0(net17),
    .A1(net9),
    .A2(net23),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG3 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[98] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.S2BEG3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG4  (.A0(net1),
    .A1(net16),
    .A2(net8),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG4 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[100] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.S2BEG4 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG5  (.A0(net2),
    .A1(net15),
    .A2(net7),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG5 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[102] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.S2BEG5 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG6  (.A0(net3),
    .A1(net14),
    .A2(net6),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG6 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[104] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.S2BEG6 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG7  (.A0(net4),
    .A1(net13),
    .A2(net5),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG7 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[106] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.S2BEG7 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG0  (.A0(net101),
    .A1(net153),
    .A2(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[2] ),
    .A3(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[3] ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[120] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W1BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG1  (.A0(net102),
    .A1(net154),
    .A2(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[3] ),
    .A3(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[2] ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[122] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W1BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG2  (.A0(net103),
    .A1(net155),
    .A2(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[0] ),
    .A3(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[1] ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[124] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W1BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG3  (.A0(net104),
    .A1(net156),
    .A2(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[1] ),
    .A3(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[0] ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[126] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W1BEG3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG0  (.A0(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[0] ),
    .A1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[0] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG0 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG7 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[128] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W2BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG1  (.A0(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[1] ),
    .A1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[1] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG1 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG6 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[130] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W2BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG2  (.A0(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[2] ),
    .A1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[2] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG2 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG5 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[132] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W2BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG3  (.A0(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[3] ),
    .A1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[3] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG3 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG4 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[134] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W2BEG3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG4  (.A0(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[0] ),
    .A1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[0] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG3 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG4 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[136] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W2BEG4 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG5  (.A0(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[1] ),
    .A1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[1] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG2 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG5 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[138] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W2BEG5 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG6  (.A0(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[2] ),
    .A1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[2] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG1 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG6 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[140] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W2BEG6 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG7  (.A0(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[3] ),
    .A1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[3] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG0 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG7 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[142] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W2BEG7 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb0  (.A0(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[0] ),
    .A1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[0] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG0 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG7 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[144] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W2BEGb0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb1  (.A0(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[1] ),
    .A1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[1] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG1 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG6 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[146] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W2BEGb1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb2  (.A0(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[2] ),
    .A1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[2] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG2 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG5 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[148] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W2BEGb2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb3  (.A0(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[3] ),
    .A1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[3] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG3 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG4 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[150] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W2BEGb3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb4  (.A0(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[0] ),
    .A1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[0] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG3 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG4 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[152] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W2BEGb4 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb5  (.A0(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[1] ),
    .A1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[1] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG2 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG5 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[154] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W2BEGb5 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb6  (.A0(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[2] ),
    .A1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[2] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG1 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG6 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[156] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W2BEGb6 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb7  (.A0(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[3] ),
    .A1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[3] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS2_BEG0 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG7 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[158] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W2BEGb7 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG0  (.A0(net121),
    .A1(net173),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG11 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG15 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[192] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[193] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W6BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG1  (.A0(net128),
    .A1(net180),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG10 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG14 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[194] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[195] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W6BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG10  (.A0(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[2] ),
    .A1(\Inst_RAM_IO_switch_matrix.J_NS4_BEG1 ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG5 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG6 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[212] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[213] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W6BEG10 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG11  (.A0(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[3] ),
    .A1(\Inst_RAM_IO_switch_matrix.J_NS4_BEG0 ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG4 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG7 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[214] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[215] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W6BEG11 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG2  (.A0(net129),
    .A1(net181),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG9 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG13 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[196] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[197] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W6BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG3  (.A0(net130),
    .A1(net182),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG8 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG12 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[198] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[199] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W6BEG3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG4  (.A0(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[0] ),
    .A1(\Inst_RAM_IO_switch_matrix.J_NS4_BEG7 ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG11 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG0 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[200] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[201] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W6BEG4 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG5  (.A0(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[1] ),
    .A1(\Inst_RAM_IO_switch_matrix.J_NS4_BEG6 ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG10 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG1 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[202] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[203] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W6BEG5 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG6  (.A0(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[2] ),
    .A1(\Inst_RAM_IO_switch_matrix.J_NS4_BEG5 ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG9 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG2 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[204] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[205] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W6BEG6 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG7  (.A0(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[3] ),
    .A1(\Inst_RAM_IO_switch_matrix.J_NS4_BEG4 ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG8 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG3 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[206] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[207] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W6BEG7 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG8  (.A0(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[0] ),
    .A1(\Inst_RAM_IO_switch_matrix.J_NS4_BEG3 ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG7 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG4 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[208] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[209] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W6BEG8 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG9  (.A0(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[1] ),
    .A1(\Inst_RAM_IO_switch_matrix.J_NS4_BEG2 ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG6 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG5 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[210] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[211] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.W6BEG9 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG0  (.A0(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[0] ),
    .A1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[0] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG15 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG7 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[160] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.WW4BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG1  (.A0(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[1] ),
    .A1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[1] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG14 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG6 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[162] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.WW4BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG10  (.A0(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[2] ),
    .A1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[2] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG5 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG5 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[180] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.WW4BEG10 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG11  (.A0(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[3] ),
    .A1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[3] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG4 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG4 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[182] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.WW4BEG11 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG12  (.A0(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[0] ),
    .A1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[0] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG3 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG3 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[184] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.WW4BEG12 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG13  (.A0(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[1] ),
    .A1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[1] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG2 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG2 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[186] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.WW4BEG13 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG14  (.A0(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[2] ),
    .A1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[2] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG1 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG1 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[188] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.WW4BEG14 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG15  (.A0(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[3] ),
    .A1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[3] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG0 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG0 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[190] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.WW4BEG15 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG2  (.A0(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[2] ),
    .A1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[2] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG13 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG5 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[164] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.WW4BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG3  (.A0(\Inst_RAM2FAB_D0_InPass4_frame_config_mux.O[3] ),
    .A1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux.O[3] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG12 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG4 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[166] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.WW4BEG3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG4  (.A0(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[0] ),
    .A1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[0] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG11 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG3 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[168] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.WW4BEG4 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG5  (.A0(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[1] ),
    .A1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[1] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG10 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG2 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[170] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.WW4BEG5 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG6  (.A0(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[2] ),
    .A1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[2] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG9 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG1 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[172] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.WW4BEG6 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG7  (.A0(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[3] ),
    .A1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[3] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG8 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG0 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[174] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.WW4BEG7 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG8  (.A0(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[0] ),
    .A1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[0] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG7 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG7 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[176] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.WW4BEG8 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG9  (.A0(\Inst_RAM2FAB_D1_InPass4_frame_config_mux.O[1] ),
    .A1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux.O[1] ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG6 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG6 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[178] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.WW4BEG9 ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._2_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._3_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.AIN[1] ),
    .B(\Inst_RAM_IO_ConfigMem.ConfigBits[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._4_  (.A1(\Inst_RAM_IO_ConfigMem.ConfigBits[74] ),
    .A2(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._0_ ),
    .B1(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.N4BEG0 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux41_buf_inst0  (.A0(net1),
    .A1(net33),
    .A2(net31),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG0 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[72] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux41_buf_inst1  (.A0(\Inst_RAM_IO_switch_matrix.J_NS4_BEG4 ),
    .A1(\Inst_RAM_IO_switch_matrix.J_NS4_BEG8 ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG12 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG0 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[72] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._2_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._3_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.AIN[1] ),
    .B(\Inst_RAM_IO_ConfigMem.ConfigBits[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._4_  (.A1(\Inst_RAM_IO_ConfigMem.ConfigBits[77] ),
    .A2(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._0_ ),
    .B1(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.N4BEG1 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux41_buf_inst0  (.A0(net2),
    .A1(net40),
    .A2(net32),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG1 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[75] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux41_buf_inst1  (.A0(\Inst_RAM_IO_switch_matrix.J_NS4_BEG5 ),
    .A1(\Inst_RAM_IO_switch_matrix.J_NS4_BEG9 ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG13 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG1 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[75] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._2_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._3_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.AIN[1] ),
    .B(\Inst_RAM_IO_ConfigMem.ConfigBits[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._4_  (.A1(\Inst_RAM_IO_ConfigMem.ConfigBits[80] ),
    .A2(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._0_ ),
    .B1(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.N4BEG2 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux41_buf_inst0  (.A0(net3),
    .A1(net41),
    .A2(net22),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG2 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[78] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux41_buf_inst1  (.A0(\Inst_RAM_IO_switch_matrix.J_NS4_BEG6 ),
    .A1(\Inst_RAM_IO_switch_matrix.J_NS4_BEG10 ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG14 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG2 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[78] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._2_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._3_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.AIN[1] ),
    .B(\Inst_RAM_IO_ConfigMem.ConfigBits[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._4_  (.A1(\Inst_RAM_IO_ConfigMem.ConfigBits[83] ),
    .A2(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._0_ ),
    .B1(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.N4BEG3 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux41_buf_inst0  (.A0(net4),
    .A1(net42),
    .A2(net23),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG3 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[81] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux41_buf_inst1  (.A0(\Inst_RAM_IO_switch_matrix.J_NS4_BEG7 ),
    .A1(\Inst_RAM_IO_switch_matrix.J_NS4_BEG11 ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG15 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG3 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[81] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._2_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._3_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.AIN[1] ),
    .B(\Inst_RAM_IO_ConfigMem.ConfigBits[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._4_  (.A1(\Inst_RAM_IO_ConfigMem.ConfigBits[110] ),
    .A2(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._0_ ),
    .B1(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.S4BEG0 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux41_buf_inst0  (.A0(net1),
    .A1(net36),
    .A2(net27),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG0 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[108] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux41_buf_inst1  (.A0(\Inst_RAM_IO_switch_matrix.J_NS4_BEG4 ),
    .A1(\Inst_RAM_IO_switch_matrix.J_NS4_BEG8 ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG12 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG4 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[108] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._2_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._3_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.AIN[1] ),
    .B(\Inst_RAM_IO_ConfigMem.ConfigBits[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._4_  (.A1(\Inst_RAM_IO_ConfigMem.ConfigBits[113] ),
    .A2(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._0_ ),
    .B1(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.S4BEG1 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux41_buf_inst0  (.A0(net2),
    .A1(net37),
    .A2(net28),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG1 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[111] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux41_buf_inst1  (.A0(\Inst_RAM_IO_switch_matrix.J_NS4_BEG5 ),
    .A1(\Inst_RAM_IO_switch_matrix.J_NS4_BEG9 ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG13 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG5 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[111] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._2_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._3_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.AIN[1] ),
    .B(\Inst_RAM_IO_ConfigMem.ConfigBits[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._4_  (.A1(\Inst_RAM_IO_ConfigMem.ConfigBits[116] ),
    .A2(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._0_ ),
    .B1(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.S4BEG2 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux41_buf_inst0  (.A0(net3),
    .A1(net38),
    .A2(net29),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG2 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[114] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux41_buf_inst1  (.A0(\Inst_RAM_IO_switch_matrix.J_NS4_BEG6 ),
    .A1(\Inst_RAM_IO_switch_matrix.J_NS4_BEG10 ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG14 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG6 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[114] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._2_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._3_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.AIN[1] ),
    .B(\Inst_RAM_IO_ConfigMem.ConfigBits[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._4_  (.A1(\Inst_RAM_IO_ConfigMem.ConfigBits[119] ),
    .A2(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._0_ ),
    .B1(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_RAM_IO_switch_matrix.S4BEG3 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux41_buf_inst0  (.A0(net4),
    .A1(net39),
    .A2(net30),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS4_BEG3 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[117] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux41_buf_inst1  (.A0(\Inst_RAM_IO_switch_matrix.J_NS4_BEG7 ),
    .A1(\Inst_RAM_IO_switch_matrix.J_NS4_BEG11 ),
    .A2(\Inst_RAM_IO_switch_matrix.J_NS4_BEG15 ),
    .A3(\Inst_RAM_IO_switch_matrix.J_NS2_BEG7 ),
    .S0(\Inst_RAM_IO_ConfigMem.ConfigBits[117] ),
    .S1(\Inst_RAM_IO_ConfigMem.ConfigBits[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_0._0_  (.A(\N4BEG_outbuf_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_0.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_1._0_  (.A(\N4BEG_outbuf_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_1.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_10._0_  (.A(\N4BEG_outbuf_10.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_10.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_11._0_  (.A(\N4BEG_outbuf_11.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_11.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_2._0_  (.A(\N4BEG_outbuf_2.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_2.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_3._0_  (.A(\N4BEG_outbuf_3.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_3.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_4._0_  (.A(\N4BEG_outbuf_4.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_5._0_  (.A(\N4BEG_outbuf_5.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_5.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_6._0_  (.A(\N4BEG_outbuf_6.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_7._0_  (.A(\N4BEG_outbuf_7.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_7.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_8._0_  (.A(\N4BEG_outbuf_8.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_8.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_9._0_  (.A(\N4BEG_outbuf_9.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_9.X ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_0._0_  (.A(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_0.A ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_1._0_  (.A(net132),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_1.A ));
 sky130_fd_sc_hd__buf_2 \N4END_inbuf_10._0_  (.A(net126),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_10.A ));
 sky130_fd_sc_hd__buf_2 \N4END_inbuf_11._0_  (.A(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_11.A ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_2._0_  (.A(net133),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_2.A ));
 sky130_fd_sc_hd__clkbuf_4 \N4END_inbuf_3._0_  (.A(net134),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_3.A ));
 sky130_fd_sc_hd__buf_2 \N4END_inbuf_4._0_  (.A(net135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_4.A ));
 sky130_fd_sc_hd__buf_2 \N4END_inbuf_5._0_  (.A(net136),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_5.A ));
 sky130_fd_sc_hd__buf_2 \N4END_inbuf_6._0_  (.A(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_6.A ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_7._0_  (.A(net123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_7.A ));
 sky130_fd_sc_hd__buf_2 \N4END_inbuf_8._0_  (.A(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_8.A ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_9._0_  (.A(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_9.A ));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__buf_2 \S4BEG_outbuf_0._0_  (.A(\S4BEG_outbuf_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_0.X ));
 sky130_fd_sc_hd__buf_2 \S4BEG_outbuf_1._0_  (.A(\S4BEG_outbuf_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_1.X ));
 sky130_fd_sc_hd__clkbuf_2 \S4BEG_outbuf_10._0_  (.A(\S4BEG_outbuf_10.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_10.X ));
 sky130_fd_sc_hd__clkbuf_2 \S4BEG_outbuf_11._0_  (.A(\S4BEG_outbuf_11.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_11.X ));
 sky130_fd_sc_hd__buf_2 \S4BEG_outbuf_2._0_  (.A(\S4BEG_outbuf_2.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_2.X ));
 sky130_fd_sc_hd__clkbuf_2 \S4BEG_outbuf_3._0_  (.A(\S4BEG_outbuf_3.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_3.X ));
 sky130_fd_sc_hd__buf_2 \S4BEG_outbuf_4._0_  (.A(\S4BEG_outbuf_4.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_2 \S4BEG_outbuf_5._0_  (.A(\S4BEG_outbuf_5.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_5.X ));
 sky130_fd_sc_hd__buf_2 \S4BEG_outbuf_6._0_  (.A(\S4BEG_outbuf_6.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_2 \S4BEG_outbuf_7._0_  (.A(\S4BEG_outbuf_7.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_7.X ));
 sky130_fd_sc_hd__buf_2 \S4BEG_outbuf_8._0_  (.A(\S4BEG_outbuf_8.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_8.X ));
 sky130_fd_sc_hd__buf_2 \S4BEG_outbuf_9._0_  (.A(\S4BEG_outbuf_9.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_9.X ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_0._0_  (.A(net183),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_0.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_1._0_  (.A(net184),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_1.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_10._0_  (.A(net178),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_10.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_11._0_  (.A(net179),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_11.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_2._0_  (.A(net185),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_2.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_3._0_  (.A(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_3.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_4._0_  (.A(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_4.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_5._0_  (.A(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_5.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_6._0_  (.A(net174),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_6.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_7._0_  (.A(net175),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_7.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_8._0_  (.A(net176),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_8.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_9._0_  (.A(net177),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_9.A ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_1 _000_ (.A(\data_outbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_1 _001_ (.A(\data_outbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_1 _002_ (.A(\data_outbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_1 _003_ (.A(\data_outbuf_3.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_1 _004_ (.A(\data_outbuf_4.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_1 _005_ (.A(\data_outbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_1 _006_ (.A(\data_outbuf_6.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_1 _007_ (.A(\data_outbuf_7.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_1 _008_ (.A(\data_outbuf_8.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_1 _009_ (.A(\data_outbuf_9.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_1 _010_ (.A(\data_outbuf_10.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_1 _011_ (.A(\data_outbuf_11.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_1 _012_ (.A(\data_outbuf_12.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_1 _013_ (.A(\data_outbuf_13.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_1 _014_ (.A(\data_outbuf_14.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_1 _015_ (.A(\data_outbuf_15.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_1 _016_ (.A(\data_outbuf_16.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_1 _017_ (.A(\data_outbuf_17.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_1 _018_ (.A(\data_outbuf_18.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_1 _019_ (.A(\data_outbuf_19.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_1 _020_ (.A(\data_outbuf_20.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_1 _021_ (.A(\data_outbuf_21.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_1 _022_ (.A(\data_outbuf_22.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_1 _023_ (.A(\data_outbuf_23.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_1 _024_ (.A(\data_outbuf_24.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_1 _025_ (.A(\data_outbuf_25.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_1 _026_ (.A(\data_outbuf_26.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_1 _027_ (.A(\data_outbuf_27.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_1 _028_ (.A(\data_outbuf_28.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_1 _029_ (.A(\data_outbuf_29.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_1 _030_ (.A(\data_outbuf_30.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_1 _031_ (.A(\data_outbuf_31.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_1 _032_ (.A(\strobe_outbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_1 _033_ (.A(\strobe_outbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_1 _034_ (.A(\strobe_outbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_1 _035_ (.A(\strobe_outbuf_3.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_1 _036_ (.A(\strobe_outbuf_4.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_1 _037_ (.A(\strobe_outbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_1 _038_ (.A(\strobe_outbuf_6.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_1 _039_ (.A(\strobe_outbuf_7.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_1 _040_ (.A(\strobe_outbuf_8.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_1 _041_ (.A(\strobe_outbuf_9.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_1 _042_ (.A(\strobe_outbuf_10.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_1 _043_ (.A(\strobe_outbuf_11.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_1 _044_ (.A(\strobe_outbuf_12.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_1 _045_ (.A(\strobe_outbuf_13.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_1 _046_ (.A(\strobe_outbuf_14.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_1 _047_ (.A(\strobe_outbuf_15.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_1 _048_ (.A(\strobe_outbuf_16.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_1 _049_ (.A(\strobe_outbuf_17.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_1 _050_ (.A(\strobe_outbuf_18.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_1 _051_ (.A(\strobe_outbuf_19.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_1 _052_ (.A(\Inst_RAM_IO_switch_matrix.N1BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_1 _053_ (.A(\Inst_RAM_IO_switch_matrix.N1BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_1 _054_ (.A(\Inst_RAM_IO_switch_matrix.N1BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_1 _055_ (.A(\Inst_RAM_IO_switch_matrix.N1BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_1 _056_ (.A(\Inst_RAM_IO_switch_matrix.N2BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_1 _057_ (.A(\Inst_RAM_IO_switch_matrix.N2BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_1 _058_ (.A(\Inst_RAM_IO_switch_matrix.N2BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_1 _059_ (.A(\Inst_RAM_IO_switch_matrix.N2BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_1 _060_ (.A(\Inst_RAM_IO_switch_matrix.N2BEG4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_1 _061_ (.A(\Inst_RAM_IO_switch_matrix.N2BEG5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_1 _062_ (.A(\Inst_RAM_IO_switch_matrix.N2BEG6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_1 _063_ (.A(\Inst_RAM_IO_switch_matrix.N2BEG7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_1 _064_ (.A(\Inst_RAM_IO_switch_matrix.N2BEGb0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_1 _065_ (.A(\Inst_RAM_IO_switch_matrix.N2BEGb1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_1 _066_ (.A(\Inst_RAM_IO_switch_matrix.N2BEGb2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_1 _067_ (.A(\Inst_RAM_IO_switch_matrix.N2BEGb3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_1 _068_ (.A(\Inst_RAM_IO_switch_matrix.N2BEGb4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_1 _069_ (.A(\Inst_RAM_IO_switch_matrix.N2BEGb5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_1 _070_ (.A(\Inst_RAM_IO_switch_matrix.N2BEGb6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_1 _071_ (.A(\Inst_RAM_IO_switch_matrix.N2BEGb7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_1 _072_ (.A(\N4BEG_outbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_1 _073_ (.A(\N4BEG_outbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_1 _074_ (.A(\N4BEG_outbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_1 _075_ (.A(\N4BEG_outbuf_3.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_1 _076_ (.A(\N4BEG_outbuf_4.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_1 _077_ (.A(\N4BEG_outbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_1 _078_ (.A(\N4BEG_outbuf_6.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_1 _079_ (.A(\N4BEG_outbuf_7.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_1 _080_ (.A(\N4BEG_outbuf_8.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_1 _081_ (.A(\N4BEG_outbuf_9.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_1 _082_ (.A(\N4BEG_outbuf_10.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_1 _083_ (.A(\N4BEG_outbuf_11.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_1 _084_ (.A(\Inst_RAM_IO_switch_matrix.N4BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_1 _085_ (.A(\Inst_RAM_IO_switch_matrix.N4BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_1 _086_ (.A(\Inst_RAM_IO_switch_matrix.N4BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_1 _087_ (.A(\Inst_RAM_IO_switch_matrix.N4BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_1 _088_ (.A(\Inst_RAM_IO_switch_matrix.S1BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_1 _089_ (.A(\Inst_RAM_IO_switch_matrix.S1BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_1 _090_ (.A(\Inst_RAM_IO_switch_matrix.S1BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_1 _091_ (.A(\Inst_RAM_IO_switch_matrix.S1BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_1 _092_ (.A(\Inst_RAM_IO_switch_matrix.S2BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_1 _093_ (.A(\Inst_RAM_IO_switch_matrix.S2BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_1 _094_ (.A(\Inst_RAM_IO_switch_matrix.S2BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_1 _095_ (.A(\Inst_RAM_IO_switch_matrix.S2BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_1 _096_ (.A(\Inst_RAM_IO_switch_matrix.S2BEG4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_1 _097_ (.A(\Inst_RAM_IO_switch_matrix.S2BEG5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net318));
 sky130_fd_sc_hd__buf_1 _098_ (.A(\Inst_RAM_IO_switch_matrix.S2BEG6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_1 _099_ (.A(\Inst_RAM_IO_switch_matrix.S2BEG7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_1 _100_ (.A(\Inst_RAM_IO_switch_matrix.S2BEGb0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_1 _101_ (.A(\Inst_RAM_IO_switch_matrix.S2BEGb1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_1 _102_ (.A(\Inst_RAM_IO_switch_matrix.S2BEGb2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_1 _103_ (.A(\Inst_RAM_IO_switch_matrix.S2BEGb3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_1 _104_ (.A(\Inst_RAM_IO_switch_matrix.S2BEGb4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_1 _105_ (.A(\Inst_RAM_IO_switch_matrix.S2BEGb5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_1 _106_ (.A(\Inst_RAM_IO_switch_matrix.S2BEGb6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_1 _107_ (.A(\Inst_RAM_IO_switch_matrix.S2BEGb7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_1 _108_ (.A(\S4BEG_outbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_1 _109_ (.A(\S4BEG_outbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_1 _110_ (.A(\S4BEG_outbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_1 _111_ (.A(\S4BEG_outbuf_3.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_1 _112_ (.A(\S4BEG_outbuf_4.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_1 _113_ (.A(\S4BEG_outbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_1 _114_ (.A(\S4BEG_outbuf_6.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_1 _115_ (.A(\S4BEG_outbuf_7.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_1 _116_ (.A(\S4BEG_outbuf_8.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_1 _117_ (.A(\S4BEG_outbuf_9.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_1 _118_ (.A(\S4BEG_outbuf_10.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_1 _119_ (.A(\S4BEG_outbuf_11.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_1 _120_ (.A(\Inst_RAM_IO_switch_matrix.S4BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_1 _121_ (.A(\Inst_RAM_IO_switch_matrix.S4BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_1 _122_ (.A(\Inst_RAM_IO_switch_matrix.S4BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_1 _123_ (.A(\Inst_RAM_IO_switch_matrix.S4BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net335));
 sky130_fd_sc_hd__buf_1 _124_ (.A(\Inst_RAM_IO_switch_matrix.W1BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_1 _125_ (.A(\Inst_RAM_IO_switch_matrix.W1BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_1 _126_ (.A(\Inst_RAM_IO_switch_matrix.W1BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net348));
 sky130_fd_sc_hd__buf_1 _127_ (.A(\Inst_RAM_IO_switch_matrix.W1BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net349));
 sky130_fd_sc_hd__buf_1 _128_ (.A(\Inst_RAM_IO_switch_matrix.W2BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_1 _129_ (.A(\Inst_RAM_IO_switch_matrix.W2BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_1 _130_ (.A(\Inst_RAM_IO_switch_matrix.W2BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_1 _131_ (.A(\Inst_RAM_IO_switch_matrix.W2BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_1 _132_ (.A(\Inst_RAM_IO_switch_matrix.W2BEG4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_1 _133_ (.A(\Inst_RAM_IO_switch_matrix.W2BEG5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_1 _134_ (.A(\Inst_RAM_IO_switch_matrix.W2BEG6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_1 _135_ (.A(\Inst_RAM_IO_switch_matrix.W2BEG7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net357));
 sky130_fd_sc_hd__buf_1 _136_ (.A(\Inst_RAM_IO_switch_matrix.W2BEGb0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_1 _137_ (.A(\Inst_RAM_IO_switch_matrix.W2BEGb1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_1 _138_ (.A(\Inst_RAM_IO_switch_matrix.W2BEGb2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_1 _139_ (.A(\Inst_RAM_IO_switch_matrix.W2BEGb3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_1 _140_ (.A(\Inst_RAM_IO_switch_matrix.W2BEGb4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_1 _141_ (.A(\Inst_RAM_IO_switch_matrix.W2BEGb5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_1 _142_ (.A(\Inst_RAM_IO_switch_matrix.W2BEGb6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_1 _143_ (.A(\Inst_RAM_IO_switch_matrix.W2BEGb7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_1 _144_ (.A(\Inst_RAM_IO_switch_matrix.W6BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net366));
 sky130_fd_sc_hd__dlymetal6s2s_1 _145_ (.A(\Inst_RAM_IO_switch_matrix.W6BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_1 _146_ (.A(\Inst_RAM_IO_switch_matrix.W6BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_1 _147_ (.A(\Inst_RAM_IO_switch_matrix.W6BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_1 _148_ (.A(\Inst_RAM_IO_switch_matrix.W6BEG4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_1 _149_ (.A(\Inst_RAM_IO_switch_matrix.W6BEG5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_1 _150_ (.A(\Inst_RAM_IO_switch_matrix.W6BEG6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_1 _151_ (.A(\Inst_RAM_IO_switch_matrix.W6BEG7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_1 _152_ (.A(\Inst_RAM_IO_switch_matrix.W6BEG8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_1 _153_ (.A(\Inst_RAM_IO_switch_matrix.W6BEG9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_1 _154_ (.A(\Inst_RAM_IO_switch_matrix.W6BEG10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_1 _155_ (.A(\Inst_RAM_IO_switch_matrix.W6BEG11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_1 _156_ (.A(\Inst_RAM_IO_switch_matrix.WW4BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_1 _157_ (.A(\Inst_RAM_IO_switch_matrix.WW4BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_1 _158_ (.A(\Inst_RAM_IO_switch_matrix.WW4BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_1 _159_ (.A(\Inst_RAM_IO_switch_matrix.WW4BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_1 _160_ (.A(\Inst_RAM_IO_switch_matrix.WW4BEG4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_1 _161_ (.A(\Inst_RAM_IO_switch_matrix.WW4BEG5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_1 _162_ (.A(\Inst_RAM_IO_switch_matrix.WW4BEG6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_1 _163_ (.A(\Inst_RAM_IO_switch_matrix.WW4BEG7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_1 _164_ (.A(\Inst_RAM_IO_switch_matrix.WW4BEG8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_1 _165_ (.A(\Inst_RAM_IO_switch_matrix.WW4BEG9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_1 _166_ (.A(\Inst_RAM_IO_switch_matrix.WW4BEG10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_1 _167_ (.A(\Inst_RAM_IO_switch_matrix.WW4BEG11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_1 _168_ (.A(\Inst_RAM_IO_switch_matrix.WW4BEG12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_1 _169_ (.A(\Inst_RAM_IO_switch_matrix.WW4BEG13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_1 _170_ (.A(\Inst_RAM_IO_switch_matrix.WW4BEG14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_1 _171_ (.A(\Inst_RAM_IO_switch_matrix.WW4BEG15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_0._0_  (.A(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_0.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_1._0_  (.A(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_1.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_10._0_  (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_10.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_11._0_  (.A(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_11.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_12._0_  (.A(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_12.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_13._0_  (.A(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_13.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_14._0_  (.A(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_14.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_15._0_  (.A(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_15.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_16._0_  (.A(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_16.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_17._0_  (.A(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_17.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_18._0_  (.A(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_18.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_19._0_  (.A(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_19.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_2._0_  (.A(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_2.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_20._0_  (.A(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_20.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_21._0_  (.A(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_21.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_22._0_  (.A(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_22.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_23._0_  (.A(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_23.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_24._0_  (.A(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_24.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_25._0_  (.A(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_25.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_26._0_  (.A(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_26.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_27._0_  (.A(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_27.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_28._0_  (.A(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_28.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_29._0_  (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_29.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_3._0_  (.A(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_3.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_30._0_  (.A(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_30.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_31._0_  (.A(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_31.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_4._0_  (.A(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_5._0_  (.A(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_5.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_6._0_  (.A(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_7._0_  (.A(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_7.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_8._0_  (.A(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_8.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_9._0_  (.A(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_9.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_0._0_  (.A(\data_inbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_0.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_1._0_  (.A(\data_inbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_1.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_10._0_  (.A(\data_inbuf_10.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_10.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_11._0_  (.A(\data_inbuf_11.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_11.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_12._0_  (.A(\data_inbuf_12.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_12.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_13._0_  (.A(\data_inbuf_13.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_13.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_14._0_  (.A(\data_inbuf_14.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_14.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_15._0_  (.A(\data_inbuf_15.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_15.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_16._0_  (.A(\data_inbuf_16.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_16.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_17._0_  (.A(\data_inbuf_17.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_17.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_18._0_  (.A(\data_inbuf_18.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_18.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_19._0_  (.A(\data_inbuf_19.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_19.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_2._0_  (.A(\data_inbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_2.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_20._0_  (.A(\data_inbuf_20.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_20.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_21._0_  (.A(\data_inbuf_21.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_21.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_22._0_  (.A(\data_inbuf_22.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_22.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_23._0_  (.A(\data_inbuf_23.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_23.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_24._0_  (.A(\data_inbuf_24.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_24.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_25._0_  (.A(\data_inbuf_25.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_25.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_26._0_  (.A(\data_inbuf_26.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_26.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_27._0_  (.A(\data_inbuf_27.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_27.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_28._0_  (.A(\data_inbuf_28.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_28.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_29._0_  (.A(\data_inbuf_29.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_29.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_3._0_  (.A(\data_inbuf_3.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_3.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_30._0_  (.A(\data_inbuf_30.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_30.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_31._0_  (.A(\data_inbuf_31.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_31.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_4._0_  (.A(\data_inbuf_4.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_5._0_  (.A(\data_inbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_5.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_6._0_  (.A(\data_inbuf_6.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_7._0_  (.A(\data_inbuf_7.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_7.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_8._0_  (.A(\data_inbuf_8.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_8.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_9._0_  (.A(\data_inbuf_9.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_9.X ));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(E1END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(E2END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__buf_8 input100 (.A(FrameStrobe[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_2 input101 (.A(N1END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_4 input102 (.A(N1END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 input103 (.A(N1END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net103));
 sky130_fd_sc_hd__buf_2 input104 (.A(N1END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net104));
 sky130_fd_sc_hd__dlymetal6s2s_1 input105 (.A(N2END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 input106 (.A(N2END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net106));
 sky130_fd_sc_hd__buf_1 input107 (.A(N2END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net107));
 sky130_fd_sc_hd__buf_2 input108 (.A(N2END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 input109 (.A(N2END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net109));
 sky130_fd_sc_hd__buf_1 input11 (.A(E2END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input110 (.A(N2END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 input111 (.A(N2END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 input112 (.A(N2END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net112));
 sky130_fd_sc_hd__buf_2 input113 (.A(N2MID[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 input114 (.A(N2MID[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net114));
 sky130_fd_sc_hd__buf_1 input115 (.A(N2MID[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 input116 (.A(N2MID[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net116));
 sky130_fd_sc_hd__buf_2 input117 (.A(N2MID[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net117));
 sky130_fd_sc_hd__buf_1 input118 (.A(N2MID[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 input119 (.A(N2MID[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net119));
 sky130_fd_sc_hd__buf_1 input12 (.A(E2END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input120 (.A(N2MID[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 input121 (.A(N4END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(N4END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(N4END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 input124 (.A(N4END[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 input125 (.A(N4END[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(N4END[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(N4END[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net127));
 sky130_fd_sc_hd__buf_2 input128 (.A(N4END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 input129 (.A(N4END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net129));
 sky130_fd_sc_hd__buf_1 input13 (.A(E2MID[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input130 (.A(N4END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 input131 (.A(N4END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(N4END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 input133 (.A(N4END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 input134 (.A(N4END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 input135 (.A(N4END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 input136 (.A(N4END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 input137 (.A(RAM2FAB_D0_I0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net137));
 sky130_fd_sc_hd__buf_1 input138 (.A(RAM2FAB_D0_I1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net138));
 sky130_fd_sc_hd__buf_1 input139 (.A(RAM2FAB_D0_I2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net139));
 sky130_fd_sc_hd__buf_1 input14 (.A(E2MID[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input140 (.A(RAM2FAB_D0_I3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net140));
 sky130_fd_sc_hd__buf_1 input141 (.A(RAM2FAB_D1_I0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net141));
 sky130_fd_sc_hd__buf_1 input142 (.A(RAM2FAB_D1_I1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net142));
 sky130_fd_sc_hd__buf_1 input143 (.A(RAM2FAB_D1_I2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net143));
 sky130_fd_sc_hd__buf_1 input144 (.A(RAM2FAB_D1_I3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net144));
 sky130_fd_sc_hd__buf_1 input145 (.A(RAM2FAB_D2_I0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 input146 (.A(RAM2FAB_D2_I1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 input147 (.A(RAM2FAB_D2_I2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net147));
 sky130_fd_sc_hd__buf_1 input148 (.A(RAM2FAB_D2_I3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 input149 (.A(RAM2FAB_D3_I0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net149));
 sky130_fd_sc_hd__buf_1 input15 (.A(E2MID[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input150 (.A(RAM2FAB_D3_I1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net150));
 sky130_fd_sc_hd__buf_1 input151 (.A(RAM2FAB_D3_I2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 input152 (.A(RAM2FAB_D3_I3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net152));
 sky130_fd_sc_hd__buf_2 input153 (.A(S1END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net153));
 sky130_fd_sc_hd__buf_2 input154 (.A(S1END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net154));
 sky130_fd_sc_hd__buf_2 input155 (.A(S1END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net155));
 sky130_fd_sc_hd__buf_2 input156 (.A(S1END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net156));
 sky130_fd_sc_hd__buf_1 input157 (.A(S2END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net157));
 sky130_fd_sc_hd__buf_1 input158 (.A(S2END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_2 input159 (.A(S2END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(E2MID[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input160 (.A(S2END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 input161 (.A(S2END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 input162 (.A(S2END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 input163 (.A(S2END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 input164 (.A(S2END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net164));
 sky130_fd_sc_hd__buf_1 input165 (.A(S2MID[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net165));
 sky130_fd_sc_hd__buf_1 input166 (.A(S2MID[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_2 input167 (.A(S2MID[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net167));
 sky130_fd_sc_hd__buf_1 input168 (.A(S2MID[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net168));
 sky130_fd_sc_hd__buf_1 input169 (.A(S2MID[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net169));
 sky130_fd_sc_hd__buf_1 input17 (.A(E2MID[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input170 (.A(S2MID[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net170));
 sky130_fd_sc_hd__buf_2 input171 (.A(S2MID[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net171));
 sky130_fd_sc_hd__buf_1 input172 (.A(S2MID[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net172));
 sky130_fd_sc_hd__buf_2 input173 (.A(S4END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 input174 (.A(S4END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 input175 (.A(S4END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 input176 (.A(S4END[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 input177 (.A(S4END[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 input178 (.A(S4END[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 input179 (.A(S4END[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(E2MID[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input180 (.A(S4END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net180));
 sky130_fd_sc_hd__buf_2 input181 (.A(S4END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net181));
 sky130_fd_sc_hd__buf_2 input182 (.A(S4END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 input183 (.A(S4END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 input184 (.A(S4END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 input185 (.A(S4END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 input186 (.A(S4END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 input187 (.A(S4END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 input188 (.A(S4END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net188));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(E2MID[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input2 (.A(E1END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input20 (.A(E2MID[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(E6END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(E6END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 sky130_fd_sc_hd__dlymetal6s2s_1 input23 (.A(E6END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(E6END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(E6END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(E6END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(E6END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__dlymetal6s2s_1 input28 (.A(E6END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(E6END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(E1END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input30 (.A(E6END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(E6END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(E6END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(EE4END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(EE4END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(EE4END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(EE4END[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(EE4END[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(EE4END[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(EE4END[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net39));
 sky130_fd_sc_hd__buf_2 input4 (.A(E1END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input40 (.A(EE4END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(EE4END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(EE4END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(EE4END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(EE4END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(EE4END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(EE4END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(EE4END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(EE4END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 input49 (.A(FrameData[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input5 (.A(E2END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input50 (.A(FrameData[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net50));
 sky130_fd_sc_hd__buf_4 input51 (.A(FrameData[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net51));
 sky130_fd_sc_hd__buf_4 input52 (.A(FrameData[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(FrameData[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_8 input54 (.A(FrameData[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 input55 (.A(FrameData[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net55));
 sky130_fd_sc_hd__buf_4 input56 (.A(FrameData[16]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net56));
 sky130_fd_sc_hd__buf_4 input57 (.A(FrameData[17]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net57));
 sky130_fd_sc_hd__buf_4 input58 (.A(FrameData[18]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net58));
 sky130_fd_sc_hd__buf_4 input59 (.A(FrameData[19]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input6 (.A(E2END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input60 (.A(FrameData[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net60));
 sky130_fd_sc_hd__buf_4 input61 (.A(FrameData[20]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net61));
 sky130_fd_sc_hd__buf_4 input62 (.A(FrameData[21]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net62));
 sky130_fd_sc_hd__buf_4 input63 (.A(FrameData[22]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net63));
 sky130_fd_sc_hd__buf_4 input64 (.A(FrameData[23]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net64));
 sky130_fd_sc_hd__buf_4 input65 (.A(FrameData[24]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net65));
 sky130_fd_sc_hd__buf_4 input66 (.A(FrameData[25]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_8 input67 (.A(FrameData[26]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net67));
 sky130_fd_sc_hd__buf_4 input68 (.A(FrameData[27]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_8 input69 (.A(FrameData[28]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net69));
 sky130_fd_sc_hd__buf_1 input7 (.A(E2END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_8 input70 (.A(FrameData[29]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_8 input71 (.A(FrameData[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net71));
 sky130_fd_sc_hd__buf_4 input72 (.A(FrameData[30]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net72));
 sky130_fd_sc_hd__buf_4 input73 (.A(FrameData[31]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net73));
 sky130_fd_sc_hd__buf_4 input74 (.A(FrameData[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net74));
 sky130_fd_sc_hd__buf_4 input75 (.A(FrameData[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net75));
 sky130_fd_sc_hd__buf_4 input76 (.A(FrameData[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net76));
 sky130_fd_sc_hd__buf_4 input77 (.A(FrameData[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net77));
 sky130_fd_sc_hd__buf_4 input78 (.A(FrameData[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net78));
 sky130_fd_sc_hd__buf_4 input79 (.A(FrameData[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net79));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(E2END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input80 (.A(FrameData[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net80));
 sky130_fd_sc_hd__buf_8 input81 (.A(FrameStrobe[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 input82 (.A(FrameStrobe[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(FrameStrobe[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(FrameStrobe[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net84));
 sky130_fd_sc_hd__buf_1 input85 (.A(FrameStrobe[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net85));
 sky130_fd_sc_hd__buf_1 input86 (.A(FrameStrobe[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(FrameStrobe[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(FrameStrobe[16]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(FrameStrobe[17]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net89));
 sky130_fd_sc_hd__buf_1 input9 (.A(E2END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input90 (.A(FrameStrobe[18]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(FrameStrobe[19]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net91));
 sky130_fd_sc_hd__buf_8 input92 (.A(FrameStrobe[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_16 input93 (.A(FrameStrobe[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net93));
 sky130_fd_sc_hd__buf_8 input94 (.A(FrameStrobe[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net94));
 sky130_fd_sc_hd__buf_8 input95 (.A(FrameStrobe[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net95));
 sky130_fd_sc_hd__buf_8 input96 (.A(FrameStrobe[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_16 input97 (.A(FrameStrobe[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net97));
 sky130_fd_sc_hd__buf_8 input98 (.A(FrameStrobe[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net98));
 sky130_fd_sc_hd__buf_8 input99 (.A(FrameStrobe[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_16 inst_clk_buf (.A(UserCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_4 output189 (.A(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Config_accessC_bit0));
 sky130_fd_sc_hd__clkbuf_4 output190 (.A(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Config_accessC_bit1));
 sky130_fd_sc_hd__clkbuf_4 output191 (.A(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Config_accessC_bit2));
 sky130_fd_sc_hd__clkbuf_4 output192 (.A(net192),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Config_accessC_bit3));
 sky130_fd_sc_hd__clkbuf_4 output193 (.A(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_A0_O0));
 sky130_fd_sc_hd__clkbuf_4 output194 (.A(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_A0_O1));
 sky130_fd_sc_hd__buf_2 output195 (.A(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_A0_O2));
 sky130_fd_sc_hd__clkbuf_4 output196 (.A(net196),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_A0_O3));
 sky130_fd_sc_hd__clkbuf_4 output197 (.A(net197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_A1_O0));
 sky130_fd_sc_hd__clkbuf_4 output198 (.A(net198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_A1_O1));
 sky130_fd_sc_hd__clkbuf_4 output199 (.A(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_A1_O2));
 sky130_fd_sc_hd__clkbuf_4 output200 (.A(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_A1_O3));
 sky130_fd_sc_hd__clkbuf_4 output201 (.A(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_C_O0));
 sky130_fd_sc_hd__clkbuf_4 output202 (.A(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_C_O1));
 sky130_fd_sc_hd__clkbuf_4 output203 (.A(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_C_O2));
 sky130_fd_sc_hd__clkbuf_4 output204 (.A(net204),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_C_O3));
 sky130_fd_sc_hd__clkbuf_4 output205 (.A(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_D0_O0));
 sky130_fd_sc_hd__clkbuf_4 output206 (.A(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_D0_O1));
 sky130_fd_sc_hd__clkbuf_4 output207 (.A(net207),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_D0_O2));
 sky130_fd_sc_hd__clkbuf_4 output208 (.A(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_D0_O3));
 sky130_fd_sc_hd__clkbuf_4 output209 (.A(net209),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_D1_O0));
 sky130_fd_sc_hd__clkbuf_4 output210 (.A(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_D1_O1));
 sky130_fd_sc_hd__clkbuf_4 output211 (.A(net211),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_D1_O2));
 sky130_fd_sc_hd__clkbuf_4 output212 (.A(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_D1_O3));
 sky130_fd_sc_hd__clkbuf_4 output213 (.A(net213),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_D2_O0));
 sky130_fd_sc_hd__clkbuf_4 output214 (.A(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_D2_O1));
 sky130_fd_sc_hd__buf_2 output215 (.A(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_D2_O2));
 sky130_fd_sc_hd__clkbuf_4 output216 (.A(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_D2_O3));
 sky130_fd_sc_hd__clkbuf_4 output217 (.A(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_D3_O0));
 sky130_fd_sc_hd__clkbuf_4 output218 (.A(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_D3_O1));
 sky130_fd_sc_hd__clkbuf_4 output219 (.A(net219),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_D3_O2));
 sky130_fd_sc_hd__clkbuf_4 output220 (.A(net220),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FAB2RAM_D3_O3));
 sky130_fd_sc_hd__clkbuf_4 output221 (.A(net221),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__clkbuf_4 output222 (.A(net222),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output223 (.A(net223),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__clkbuf_4 output224 (.A(net224),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output225 (.A(net225),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__clkbuf_4 output226 (.A(net226),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__clkbuf_4 output227 (.A(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__clkbuf_4 output228 (.A(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__clkbuf_4 output229 (.A(net229),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__clkbuf_4 output230 (.A(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__clkbuf_4 output231 (.A(net231),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__clkbuf_4 output232 (.A(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__clkbuf_4 output233 (.A(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__clkbuf_4 output234 (.A(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__clkbuf_4 output235 (.A(net235),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__clkbuf_4 output236 (.A(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__clkbuf_4 output237 (.A(net237),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__clkbuf_4 output238 (.A(net238),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__clkbuf_4 output239 (.A(net239),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__clkbuf_4 output240 (.A(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__clkbuf_4 output241 (.A(net241),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__clkbuf_4 output242 (.A(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__clkbuf_4 output243 (.A(net243),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__clkbuf_4 output244 (.A(net244),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__clkbuf_4 output245 (.A(net245),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output246 (.A(net246),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__clkbuf_4 output247 (.A(net247),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__clkbuf_4 output248 (.A(net248),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__clkbuf_4 output249 (.A(net249),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__clkbuf_4 output250 (.A(net250),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__clkbuf_4 output251 (.A(net251),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__clkbuf_4 output252 (.A(net252),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output253 (.A(net253),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__clkbuf_4 output254 (.A(net254),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__clkbuf_4 output255 (.A(net255),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__clkbuf_4 output256 (.A(net256),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__clkbuf_4 output257 (.A(net257),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__clkbuf_4 output258 (.A(net258),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__clkbuf_4 output259 (.A(net259),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__clkbuf_4 output260 (.A(net260),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__clkbuf_4 output261 (.A(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__clkbuf_4 output262 (.A(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__clkbuf_4 output263 (.A(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__clkbuf_4 output264 (.A(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__clkbuf_4 output265 (.A(net265),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__clkbuf_4 output266 (.A(net266),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__buf_2 output267 (.A(net267),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__clkbuf_4 output268 (.A(net268),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__buf_2 output269 (.A(net269),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__clkbuf_4 output270 (.A(net270),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__clkbuf_4 output271 (.A(net271),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__clkbuf_4 output272 (.A(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_2 output273 (.A(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output274 (.A(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output275 (.A(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output276 (.A(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output277 (.A(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output278 (.A(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output279 (.A(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output280 (.A(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEG[3]));
 sky130_fd_sc_hd__buf_2 output281 (.A(net281),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEG[4]));
 sky130_fd_sc_hd__buf_2 output282 (.A(net282),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output283 (.A(net283),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output284 (.A(net284),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output285 (.A(net285),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output286 (.A(net286),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEGb[1]));
 sky130_fd_sc_hd__clkbuf_4 output287 (.A(net287),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output288 (.A(net288),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEGb[3]));
 sky130_fd_sc_hd__clkbuf_4 output289 (.A(net289),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output290 (.A(net290),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEGb[5]));
 sky130_fd_sc_hd__clkbuf_4 output291 (.A(net291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEGb[6]));
 sky130_fd_sc_hd__clkbuf_4 output292 (.A(net292),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEGb[7]));
 sky130_fd_sc_hd__clkbuf_4 output293 (.A(net293),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output294 (.A(net294),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[10]));
 sky130_fd_sc_hd__buf_2 output295 (.A(net295),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output296 (.A(net296),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output297 (.A(net297),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output298 (.A(net298),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output299 (.A(net299),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[15]));
 sky130_fd_sc_hd__buf_2 output300 (.A(net300),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output301 (.A(net301),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[2]));
 sky130_fd_sc_hd__buf_2 output302 (.A(net302),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output303 (.A(net303),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output304 (.A(net304),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output305 (.A(net305),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output306 (.A(net306),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output307 (.A(net307),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[8]));
 sky130_fd_sc_hd__buf_2 output308 (.A(net308),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output309 (.A(net309),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S1BEG[0]));
 sky130_fd_sc_hd__buf_2 output310 (.A(net310),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output311 (.A(net311),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output312 (.A(net312),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output313 (.A(net313),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEG[0]));
 sky130_fd_sc_hd__buf_2 output314 (.A(net314),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output315 (.A(net315),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEG[2]));
 sky130_fd_sc_hd__buf_2 output316 (.A(net316),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEG[3]));
 sky130_fd_sc_hd__buf_2 output317 (.A(net317),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output318 (.A(net318),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output319 (.A(net319),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEG[6]));
 sky130_fd_sc_hd__buf_2 output320 (.A(net320),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output321 (.A(net321),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output322 (.A(net322),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEGb[1]));
 sky130_fd_sc_hd__clkbuf_4 output323 (.A(net323),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output324 (.A(net324),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEGb[3]));
 sky130_fd_sc_hd__clkbuf_4 output325 (.A(net325),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output326 (.A(net326),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEGb[5]));
 sky130_fd_sc_hd__clkbuf_4 output327 (.A(net327),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEGb[6]));
 sky130_fd_sc_hd__clkbuf_4 output328 (.A(net328),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output329 (.A(net329),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output330 (.A(net330),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output331 (.A(net331),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output332 (.A(net332),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output333 (.A(net333),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output334 (.A(net334),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output335 (.A(net335),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output336 (.A(net336),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output337 (.A(net337),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output338 (.A(net338),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output339 (.A(net339),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output340 (.A(net340),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output341 (.A(net341),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[6]));
 sky130_fd_sc_hd__buf_2 output342 (.A(net342),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output343 (.A(net343),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output344 (.A(net344),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[9]));
 sky130_fd_sc_hd__buf_1 output345 (.A(net345),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(UserCLKo));
 sky130_fd_sc_hd__clkbuf_4 output346 (.A(net346),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output347 (.A(net347),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output348 (.A(net348),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output349 (.A(net349),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output350 (.A(net350),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output351 (.A(net351),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output352 (.A(net352),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output353 (.A(net353),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output354 (.A(net354),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output355 (.A(net355),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output356 (.A(net356),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output357 (.A(net357),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output358 (.A(net358),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output359 (.A(net359),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEGb[1]));
 sky130_fd_sc_hd__clkbuf_4 output360 (.A(net360),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEGb[2]));
 sky130_fd_sc_hd__clkbuf_4 output361 (.A(net361),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEGb[3]));
 sky130_fd_sc_hd__clkbuf_4 output362 (.A(net362),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output363 (.A(net363),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEGb[5]));
 sky130_fd_sc_hd__clkbuf_4 output364 (.A(net364),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEGb[6]));
 sky130_fd_sc_hd__clkbuf_4 output365 (.A(net365),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEGb[7]));
 sky130_fd_sc_hd__clkbuf_4 output366 (.A(net366),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output367 (.A(net367),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output368 (.A(net368),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output369 (.A(net369),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output370 (.A(net370),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output371 (.A(net371),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output372 (.A(net372),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output373 (.A(net373),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output374 (.A(net374),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output375 (.A(net375),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output376 (.A(net376),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output377 (.A(net377),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output378 (.A(net378),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output379 (.A(net379),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output380 (.A(net380),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output381 (.A(net381),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output382 (.A(net382),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output383 (.A(net383),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output384 (.A(net384),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output385 (.A(net385),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output386 (.A(net386),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output387 (.A(net387),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output388 (.A(net388),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output389 (.A(net389),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output390 (.A(net390),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output391 (.A(net391),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output392 (.A(net392),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output393 (.A(net393),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[9]));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_0._0_  (.A(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_0.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_1._0_  (.A(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_1.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_10._0_  (.A(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_10.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_11._0_  (.A(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_11.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_12._0_  (.A(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_12.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_13._0_  (.A(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_13.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_14._0_  (.A(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_14.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_15._0_  (.A(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_15.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_16._0_  (.A(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_16.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_17._0_  (.A(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_17.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_18._0_  (.A(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_18.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_19._0_  (.A(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_19.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_2._0_  (.A(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_2.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_3._0_  (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_3.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_4._0_  (.A(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_5._0_  (.A(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_5.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_6._0_  (.A(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_7._0_  (.A(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_7.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_8._0_  (.A(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_8.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_9._0_  (.A(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_9.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_0._0_  (.A(\strobe_inbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_0.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_1._0_  (.A(\strobe_inbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_1.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_10._0_  (.A(\strobe_inbuf_10.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_10.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_11._0_  (.A(\strobe_inbuf_11.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_11.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_12._0_  (.A(\strobe_inbuf_12.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_12.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_13._0_  (.A(\strobe_inbuf_13.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_13.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_14._0_  (.A(\strobe_inbuf_14.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_14.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_15._0_  (.A(\strobe_inbuf_15.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_15.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_16._0_  (.A(\strobe_inbuf_16.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_16.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_17._0_  (.A(\strobe_inbuf_17.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_17.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_18._0_  (.A(\strobe_inbuf_18.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_18.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_19._0_  (.A(\strobe_inbuf_19.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_19.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_2._0_  (.A(\strobe_inbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_2.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_3._0_  (.A(\strobe_inbuf_3.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_3.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_4._0_  (.A(\strobe_inbuf_4.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_5._0_  (.A(\strobe_inbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_5.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_6._0_  (.A(\strobe_inbuf_6.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_7._0_  (.A(\strobe_inbuf_7.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_7.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_8._0_  (.A(\strobe_inbuf_8.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_8.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_9._0_  (.A(\strobe_inbuf_9.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_9.X ));
endmodule
