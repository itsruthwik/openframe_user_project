module N_term_single2 (UserCLK,
    UserCLKo,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1END,
    N2END,
    N2MID,
    N4END,
    NN4END,
    S1BEG,
    S2BEG,
    S2BEGb,
    S4BEG,
    SS4BEG);
 input UserCLK;
 output UserCLKo;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 input [3:0] N1END;
 input [7:0] N2END;
 input [7:0] N2MID;
 input [15:0] N4END;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 output [15:0] S4BEG;
 output [15:0] SS4BEG;

 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;

 sky130_fd_sc_hd__clkbuf_2 _000_ (.A(FrameData[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 _001_ (.A(FrameData[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 _002_ (.A(FrameData[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 _003_ (.A(FrameData[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 _004_ (.A(FrameData[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 _005_ (.A(FrameData[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 _006_ (.A(FrameData[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 _007_ (.A(FrameData[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 _008_ (.A(FrameData[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 _009_ (.A(FrameData[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 _010_ (.A(FrameData[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 _011_ (.A(FrameData[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 _012_ (.A(FrameData[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 _013_ (.A(FrameData[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 _014_ (.A(FrameData[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 _015_ (.A(FrameData[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 _016_ (.A(FrameData[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 _017_ (.A(FrameData[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 _018_ (.A(FrameData[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 _019_ (.A(FrameData[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 _020_ (.A(FrameData[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 _021_ (.A(FrameData[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 _022_ (.A(FrameData[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 _023_ (.A(FrameData[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 _024_ (.A(FrameData[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 _025_ (.A(FrameData[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 _026_ (.A(FrameData[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 _027_ (.A(FrameData[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 _028_ (.A(FrameData[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 _029_ (.A(FrameData[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 _030_ (.A(FrameData[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 _031_ (.A(FrameData[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 _032_ (.A(FrameStrobe[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 _033_ (.A(FrameStrobe[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 _034_ (.A(FrameStrobe[2]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 _035_ (.A(FrameStrobe[3]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 _036_ (.A(FrameStrobe[4]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 _037_ (.A(FrameStrobe[5]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 _038_ (.A(FrameStrobe[6]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 _039_ (.A(FrameStrobe[7]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 _040_ (.A(FrameStrobe[8]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 _041_ (.A(FrameStrobe[9]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 _042_ (.A(FrameStrobe[10]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 _043_ (.A(FrameStrobe[11]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 _044_ (.A(FrameStrobe[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 _045_ (.A(FrameStrobe[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 _046_ (.A(FrameStrobe[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 _047_ (.A(FrameStrobe[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 _048_ (.A(FrameStrobe[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 _049_ (.A(FrameStrobe[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 _050_ (.A(FrameStrobe[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 _051_ (.A(FrameStrobe[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 _052_ (.A(N1END[3]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 _053_ (.A(N1END[2]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 _054_ (.A(N1END[1]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 _055_ (.A(N1END[0]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 _056_ (.A(N2MID[7]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 _057_ (.A(N2MID[6]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 _058_ (.A(N2MID[5]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 _059_ (.A(N2MID[4]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 _060_ (.A(N2MID[3]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 _061_ (.A(N2MID[2]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 _062_ (.A(N2MID[1]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 _063_ (.A(N2MID[0]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 _064_ (.A(N2END[7]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 _065_ (.A(N2END[6]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 _066_ (.A(N2END[5]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 _067_ (.A(N2END[4]),
    .X(net68));
 sky130_fd_sc_hd__buf_1 _068_ (.A(N2END[3]),
    .X(net69));
 sky130_fd_sc_hd__buf_1 _069_ (.A(N2END[2]),
    .X(net70));
 sky130_fd_sc_hd__buf_1 _070_ (.A(N2END[1]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 _071_ (.A(N2END[0]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 _072_ (.A(N4END[15]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 _073_ (.A(N4END[14]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _074_ (.A(N4END[13]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 _075_ (.A(N4END[12]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 _076_ (.A(N4END[11]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 _077_ (.A(N4END[10]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 _078_ (.A(N4END[9]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 _079_ (.A(N4END[8]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 _080_ (.A(N4END[7]),
    .X(net87));
 sky130_fd_sc_hd__buf_1 _081_ (.A(N4END[6]),
    .X(net88));
 sky130_fd_sc_hd__buf_1 _082_ (.A(N4END[5]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 _083_ (.A(N4END[4]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 _084_ (.A(N4END[3]),
    .X(net76));
 sky130_fd_sc_hd__buf_1 _085_ (.A(N4END[2]),
    .X(net77));
 sky130_fd_sc_hd__buf_1 _086_ (.A(N4END[1]),
    .X(net78));
 sky130_fd_sc_hd__buf_1 _087_ (.A(N4END[0]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 _088_ (.A(NN4END[15]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 _089_ (.A(NN4END[14]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 _090_ (.A(NN4END[13]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 _091_ (.A(NN4END[12]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 _092_ (.A(NN4END[11]),
    .X(net99));
 sky130_fd_sc_hd__buf_1 _093_ (.A(NN4END[10]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 _094_ (.A(NN4END[9]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 _095_ (.A(NN4END[8]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 _096_ (.A(NN4END[7]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 _097_ (.A(NN4END[6]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 _098_ (.A(NN4END[5]),
    .X(net90));
 sky130_fd_sc_hd__buf_1 _099_ (.A(NN4END[4]),
    .X(net91));
 sky130_fd_sc_hd__buf_1 _100_ (.A(NN4END[3]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 _101_ (.A(NN4END[2]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 _102_ (.A(NN4END[1]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 _103_ (.A(NN4END[0]),
    .X(net95));
 sky130_fd_sc_hd__buf_2 _104_ (.A(UserCLK),
    .X(net105));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_135 ();
 sky130_fd_sc_hd__buf_2 output1 (.A(net1),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output2 (.A(net2),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output3 (.A(net3),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(S1BEG[0]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(S1BEG[1]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(S1BEG[2]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(S1BEG[3]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(S2BEG[0]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(S2BEG[1]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(S2BEG[2]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(S2BEG[3]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(S2BEG[4]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(S2BEG[5]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(S2BEG[6]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(S2BEG[7]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(S2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(S2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(S2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(S2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(S2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(S2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(S2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(S2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(S4BEG[0]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(S4BEG[10]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(S4BEG[11]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(S4BEG[12]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(S4BEG[13]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(S4BEG[14]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(S4BEG[15]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(S4BEG[1]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(S4BEG[2]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(S4BEG[3]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(S4BEG[4]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(S4BEG[5]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(S4BEG[6]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(S4BEG[7]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(S4BEG[8]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(S4BEG[9]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(SS4BEG[0]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(SS4BEG[10]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(SS4BEG[11]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(SS4BEG[12]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(SS4BEG[13]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(SS4BEG[14]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(SS4BEG[15]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(SS4BEG[1]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(SS4BEG[2]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(SS4BEG[3]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(SS4BEG[4]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(SS4BEG[5]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(SS4BEG[6]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(SS4BEG[7]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(SS4BEG[8]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(SS4BEG[9]));
 sky130_fd_sc_hd__buf_1 output105 (.A(net105),
    .X(UserCLKo));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(FrameData[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(FrameData[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(FrameData[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(FrameData[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(FrameData[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(FrameData[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(FrameData[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(FrameData[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(FrameData[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(FrameData[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(FrameData[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(FrameData[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(FrameData[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(FrameData[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(FrameStrobe[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(N4END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(N4END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(N4END[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(N4END[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(N4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(NN4END[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(NN4END[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(NN4END[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(NN4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(N2END[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(NN4END[11]));
 sky130_fd_sc_hd__decap_3 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_472 ();
endmodule
