magic
tech sky130A
magscale 1 2
timestamp 1746770486
<< viali >>
rect 1593 8585 1627 8619
rect 3249 8585 3283 8619
rect 4813 8585 4847 8619
rect 6469 8585 6503 8619
rect 7941 8585 7975 8619
rect 9505 8585 9539 8619
rect 12633 8585 12667 8619
rect 14197 8585 14231 8619
rect 15761 8585 15795 8619
rect 17325 8585 17359 8619
rect 18889 8585 18923 8619
rect 20453 8585 20487 8619
rect 22017 8585 22051 8619
rect 23581 8585 23615 8619
rect 25237 8585 25271 8619
rect 27077 8585 27111 8619
rect 28273 8585 28307 8619
rect 29929 8585 29963 8619
rect 31125 8585 31159 8619
rect 31493 8585 31527 8619
rect 32873 8585 32907 8619
rect 1777 8449 1811 8483
rect 3433 8449 3467 8483
rect 4997 8449 5031 8483
rect 6653 8449 6687 8483
rect 8125 8449 8159 8483
rect 9689 8449 9723 8483
rect 11253 8449 11287 8483
rect 12817 8449 12851 8483
rect 14381 8449 14415 8483
rect 15945 8449 15979 8483
rect 17509 8449 17543 8483
rect 19073 8449 19107 8483
rect 20637 8449 20671 8483
rect 22201 8449 22235 8483
rect 23765 8449 23799 8483
rect 25053 8449 25087 8483
rect 27261 8449 27295 8483
rect 28457 8449 28491 8483
rect 29745 8449 29779 8483
rect 30941 8449 30975 8483
rect 31309 8449 31343 8483
rect 31677 8449 31711 8483
rect 32321 8449 32355 8483
rect 32689 8449 32723 8483
rect 11069 8313 11103 8347
rect 31861 8313 31895 8347
rect 32505 8245 32539 8279
rect 31401 8041 31435 8075
rect 31769 8041 31803 8075
rect 32137 8041 32171 8075
rect 31217 7837 31251 7871
rect 31585 7837 31619 7871
rect 31953 7837 31987 7871
rect 32321 7837 32355 7871
rect 32689 7837 32723 7871
rect 32505 7701 32539 7735
rect 32873 7701 32907 7735
rect 9321 7497 9355 7531
rect 11069 7497 11103 7531
rect 14197 7497 14231 7531
rect 14841 7497 14875 7531
rect 17601 7497 17635 7531
rect 19993 7497 20027 7531
rect 24409 7497 24443 7531
rect 24777 7497 24811 7531
rect 25329 7497 25363 7531
rect 27721 7497 27755 7531
rect 27997 7497 28031 7531
rect 28273 7497 28307 7531
rect 28549 7497 28583 7531
rect 29469 7497 29503 7531
rect 30941 7497 30975 7531
rect 32505 7497 32539 7531
rect 9229 7361 9263 7395
rect 9505 7361 9539 7395
rect 11253 7361 11287 7395
rect 12357 7361 12391 7395
rect 14381 7361 14415 7395
rect 14749 7361 14783 7395
rect 15025 7361 15059 7395
rect 17693 7361 17727 7395
rect 17785 7361 17819 7395
rect 18061 7361 18095 7395
rect 19809 7361 19843 7395
rect 21833 7361 21867 7395
rect 22385 7361 22419 7395
rect 22477 7361 22511 7395
rect 23949 7361 23983 7395
rect 24225 7361 24259 7395
rect 24501 7361 24535 7395
rect 24961 7361 24995 7395
rect 25513 7361 25547 7395
rect 27905 7361 27939 7395
rect 28181 7361 28215 7395
rect 28457 7361 28491 7395
rect 28733 7361 28767 7395
rect 29653 7361 29687 7395
rect 31125 7361 31159 7395
rect 32321 7361 32355 7395
rect 32689 7361 32723 7395
rect 10885 7293 10919 7327
rect 24685 7225 24719 7259
rect 12173 7157 12207 7191
rect 17969 7157 18003 7191
rect 18245 7157 18279 7191
rect 22017 7157 22051 7191
rect 22293 7157 22327 7191
rect 22661 7157 22695 7191
rect 24133 7157 24167 7191
rect 32873 7157 32907 7191
rect 21649 6885 21683 6919
rect 20729 6817 20763 6851
rect 20269 6749 20303 6783
rect 21097 6749 21131 6783
rect 21189 6749 21223 6783
rect 21465 6749 21499 6783
rect 24593 6749 24627 6783
rect 24685 6749 24719 6783
rect 25329 6749 25363 6783
rect 26249 6749 26283 6783
rect 28917 6749 28951 6783
rect 32321 6749 32355 6783
rect 32689 6749 32723 6783
rect 21005 6681 21039 6715
rect 20453 6613 20487 6647
rect 21373 6613 21407 6647
rect 24409 6613 24443 6647
rect 24869 6613 24903 6647
rect 25145 6613 25179 6647
rect 26065 6613 26099 6647
rect 28733 6613 28767 6647
rect 32505 6613 32539 6647
rect 32873 6613 32907 6647
rect 19165 6409 19199 6443
rect 29745 6409 29779 6443
rect 32873 6409 32907 6443
rect 18521 6341 18555 6375
rect 18153 6273 18187 6307
rect 18705 6273 18739 6307
rect 18981 6273 19015 6307
rect 29929 6273 29963 6307
rect 32321 6273 32355 6307
rect 32689 6273 32723 6307
rect 18613 6137 18647 6171
rect 18889 6137 18923 6171
rect 18337 6069 18371 6103
rect 19257 6069 19291 6103
rect 32505 6069 32539 6103
rect 17049 5865 17083 5899
rect 31033 5865 31067 5899
rect 32873 5797 32907 5831
rect 17785 5729 17819 5763
rect 17141 5661 17175 5695
rect 17233 5661 17267 5695
rect 17509 5661 17543 5695
rect 30849 5661 30883 5695
rect 32321 5661 32355 5695
rect 32689 5661 32723 5695
rect 17417 5525 17451 5559
rect 17693 5525 17727 5559
rect 32505 5525 32539 5559
rect 15577 5321 15611 5355
rect 16405 5321 16439 5355
rect 16957 5321 16991 5355
rect 32873 5321 32907 5355
rect 15301 5185 15335 5219
rect 15393 5185 15427 5219
rect 16497 5185 16531 5219
rect 16773 5185 16807 5219
rect 17049 5185 17083 5219
rect 17325 5185 17359 5219
rect 28733 5185 28767 5219
rect 32321 5185 32355 5219
rect 32689 5185 32723 5219
rect 17233 5049 17267 5083
rect 28917 5049 28951 5083
rect 32505 4981 32539 5015
rect 3157 4777 3191 4811
rect 3433 4777 3467 4811
rect 7389 4777 7423 4811
rect 12081 4777 12115 4811
rect 13553 4777 13587 4811
rect 15393 4777 15427 4811
rect 15945 4777 15979 4811
rect 16221 4777 16255 4811
rect 13277 4709 13311 4743
rect 15209 4709 15243 4743
rect 16589 4709 16623 4743
rect 28733 4709 28767 4743
rect 32873 4709 32907 4743
rect 2973 4573 3007 4607
rect 3249 4573 3283 4607
rect 3801 4573 3835 4607
rect 7205 4573 7239 4607
rect 10793 4573 10827 4607
rect 11069 4573 11103 4607
rect 11345 4573 11379 4607
rect 11621 4573 11655 4607
rect 11897 4573 11931 4607
rect 12265 4573 12299 4607
rect 12541 4573 12575 4607
rect 13093 4573 13127 4607
rect 13369 4573 13403 4607
rect 13645 4573 13679 4607
rect 14749 4573 14783 4607
rect 15025 4573 15059 4607
rect 15393 4573 15427 4607
rect 15485 4573 15519 4607
rect 15761 4573 15795 4607
rect 16037 4573 16071 4607
rect 16313 4573 16347 4607
rect 16405 4573 16439 4607
rect 27905 4573 27939 4607
rect 28273 4573 28307 4607
rect 28641 4573 28675 4607
rect 28917 4573 28951 4607
rect 32321 4573 32355 4607
rect 32689 4573 32723 4607
rect 27997 4505 28031 4539
rect 3985 4437 4019 4471
rect 10977 4437 11011 4471
rect 11253 4437 11287 4471
rect 11529 4437 11563 4471
rect 11805 4437 11839 4471
rect 12449 4437 12483 4471
rect 12725 4437 12759 4471
rect 13829 4437 13863 4471
rect 14933 4437 14967 4471
rect 15669 4437 15703 4471
rect 27721 4437 27755 4471
rect 28457 4437 28491 4471
rect 32505 4437 32539 4471
rect 2697 4233 2731 4267
rect 3157 4233 3191 4267
rect 7021 4233 7055 4267
rect 29377 4233 29411 4267
rect 1961 4097 1995 4131
rect 2237 4097 2271 4131
rect 2513 4097 2547 4131
rect 2973 4097 3007 4131
rect 3433 4097 3467 4131
rect 3709 4097 3743 4131
rect 4261 4097 4295 4131
rect 4629 4097 4663 4131
rect 6561 4097 6595 4131
rect 6837 4097 6871 4131
rect 7113 4097 7147 4131
rect 7389 4097 7423 4131
rect 7665 4097 7699 4131
rect 7941 4097 7975 4131
rect 14013 4097 14047 4131
rect 14473 4097 14507 4131
rect 15117 4097 15151 4131
rect 15393 4097 15427 4131
rect 27169 4097 27203 4131
rect 27537 4097 27571 4131
rect 27721 4097 27755 4131
rect 27997 4097 28031 4131
rect 28273 4097 28307 4131
rect 28549 4097 28583 4131
rect 28825 4097 28859 4131
rect 29101 4097 29135 4131
rect 29193 4097 29227 4131
rect 29561 4097 29595 4131
rect 32321 4097 32355 4131
rect 32689 4097 32723 4131
rect 28457 4029 28491 4063
rect 2421 3961 2455 3995
rect 4813 3961 4847 3995
rect 15577 3961 15611 3995
rect 28089 3961 28123 3995
rect 32873 3961 32907 3995
rect 2145 3893 2179 3927
rect 3617 3893 3651 3927
rect 3893 3893 3927 3927
rect 4445 3893 4479 3927
rect 6745 3893 6779 3927
rect 7297 3893 7331 3927
rect 7573 3893 7607 3927
rect 7849 3893 7883 3927
rect 8125 3893 8159 3927
rect 14197 3893 14231 3927
rect 14657 3893 14691 3927
rect 15301 3893 15335 3927
rect 26985 3893 27019 3927
rect 27537 3893 27571 3927
rect 27813 3893 27847 3927
rect 28641 3893 28675 3927
rect 28917 3893 28951 3927
rect 29193 3893 29227 3927
rect 32505 3893 32539 3927
rect 23765 3689 23799 3723
rect 24133 3689 24167 3723
rect 24869 3689 24903 3723
rect 19441 3621 19475 3655
rect 21189 3621 21223 3655
rect 21465 3621 21499 3655
rect 25145 3621 25179 3655
rect 32873 3621 32907 3655
rect 20729 3553 20763 3587
rect 25237 3553 25271 3587
rect 2329 3485 2363 3519
rect 7205 3485 7239 3519
rect 17877 3485 17911 3519
rect 17969 3485 18003 3519
rect 19257 3485 19291 3519
rect 20913 3485 20947 3519
rect 21005 3485 21039 3519
rect 21281 3485 21315 3519
rect 21566 3485 21600 3519
rect 21833 3485 21867 3519
rect 22293 3485 22327 3519
rect 23673 3485 23707 3519
rect 23949 3485 23983 3519
rect 24409 3485 24443 3519
rect 24685 3485 24719 3519
rect 24961 3485 24995 3519
rect 25421 3485 25455 3519
rect 26617 3485 26651 3519
rect 26893 3485 26927 3519
rect 27445 3485 27479 3519
rect 27721 3485 27755 3519
rect 28181 3485 28215 3519
rect 28457 3485 28491 3519
rect 28549 3485 28583 3519
rect 32321 3485 32355 3519
rect 32689 3485 32723 3519
rect 19533 3417 19567 3451
rect 23857 3417 23891 3451
rect 27813 3417 27847 3451
rect 2513 3349 2547 3383
rect 7389 3349 7423 3383
rect 17785 3349 17819 3383
rect 18153 3349 18187 3383
rect 20821 3349 20855 3383
rect 21741 3349 21775 3383
rect 22017 3349 22051 3383
rect 22201 3349 22235 3383
rect 23581 3349 23615 3383
rect 24593 3349 24627 3383
rect 26433 3349 26467 3383
rect 26709 3349 26743 3383
rect 27261 3349 27295 3383
rect 27537 3349 27571 3383
rect 27997 3349 28031 3383
rect 28273 3349 28307 3383
rect 28549 3349 28583 3383
rect 32505 3349 32539 3383
rect 22661 3145 22695 3179
rect 24501 3145 24535 3179
rect 25605 3145 25639 3179
rect 27629 3145 27663 3179
rect 32873 3145 32907 3179
rect 15485 3009 15519 3043
rect 15853 3009 15887 3043
rect 16221 3009 16255 3043
rect 16773 3009 16807 3043
rect 17141 3009 17175 3043
rect 17509 3009 17543 3043
rect 18981 3009 19015 3043
rect 19349 3009 19383 3043
rect 19717 3009 19751 3043
rect 20085 3009 20119 3043
rect 20453 3009 20487 3043
rect 20821 3009 20855 3043
rect 21189 3009 21223 3043
rect 21833 3009 21867 3043
rect 22201 3009 22235 3043
rect 22845 3009 22879 3043
rect 23213 3009 23247 3043
rect 23581 3009 23615 3043
rect 23949 3009 23983 3043
rect 24317 3009 24351 3043
rect 24685 3009 24719 3043
rect 25053 3009 25087 3043
rect 25421 3009 25455 3043
rect 25789 3009 25823 3043
rect 27813 3009 27847 3043
rect 31677 3009 31711 3043
rect 32321 3009 32355 3043
rect 32689 3009 32723 3043
rect 20269 2873 20303 2907
rect 21005 2873 21039 2907
rect 22385 2873 22419 2907
rect 23029 2873 23063 2907
rect 23765 2873 23799 2907
rect 24869 2873 24903 2907
rect 25237 2873 25271 2907
rect 15669 2805 15703 2839
rect 16037 2805 16071 2839
rect 16405 2805 16439 2839
rect 16957 2805 16991 2839
rect 17325 2805 17359 2839
rect 17693 2805 17727 2839
rect 19165 2805 19199 2839
rect 19533 2805 19567 2839
rect 19901 2805 19935 2839
rect 20637 2805 20671 2839
rect 21373 2805 21407 2839
rect 22017 2805 22051 2839
rect 23397 2805 23431 2839
rect 24133 2805 24167 2839
rect 31861 2805 31895 2839
rect 32505 2805 32539 2839
rect 19441 2601 19475 2635
rect 21281 2601 21315 2635
rect 23765 2601 23799 2635
rect 25605 2601 25639 2635
rect 14933 2533 14967 2567
rect 16037 2533 16071 2567
rect 18981 2533 19015 2567
rect 20545 2533 20579 2567
rect 22017 2533 22051 2567
rect 23397 2533 23431 2567
rect 24869 2533 24903 2567
rect 25237 2533 25271 2567
rect 32873 2533 32907 2567
rect 14749 2397 14783 2431
rect 15117 2397 15151 2431
rect 15485 2397 15519 2431
rect 15853 2397 15887 2431
rect 16221 2397 16255 2431
rect 16957 2397 16991 2431
rect 17325 2397 17359 2431
rect 17693 2397 17727 2431
rect 18061 2397 18095 2431
rect 18429 2397 18463 2431
rect 18797 2397 18831 2431
rect 19257 2397 19291 2431
rect 19625 2397 19659 2431
rect 19993 2397 20027 2431
rect 20361 2397 20395 2431
rect 20729 2397 20763 2431
rect 21097 2397 21131 2431
rect 21833 2397 21867 2431
rect 22201 2397 22235 2431
rect 22569 2397 22603 2431
rect 22937 2397 22971 2431
rect 23581 2397 23615 2431
rect 23949 2397 23983 2431
rect 24685 2397 24719 2431
rect 25053 2397 25087 2431
rect 25421 2397 25455 2431
rect 25789 2397 25823 2431
rect 26157 2397 26191 2431
rect 30941 2397 30975 2431
rect 31309 2397 31343 2431
rect 31677 2397 31711 2431
rect 32321 2397 32355 2431
rect 32689 2397 32723 2431
rect 15301 2261 15335 2295
rect 15669 2261 15703 2295
rect 16405 2261 16439 2295
rect 17141 2261 17175 2295
rect 17509 2261 17543 2295
rect 17877 2261 17911 2295
rect 18245 2261 18279 2295
rect 18613 2261 18647 2295
rect 19809 2261 19843 2295
rect 20177 2261 20211 2295
rect 20913 2261 20947 2295
rect 22385 2261 22419 2295
rect 22753 2261 22787 2295
rect 23121 2261 23155 2295
rect 24501 2261 24535 2295
rect 25973 2261 26007 2295
rect 31125 2261 31159 2295
rect 31493 2261 31527 2295
rect 31861 2261 31895 2295
rect 32505 2261 32539 2295
<< metal1 >>
rect 14366 9052 14372 9104
rect 14424 9092 14430 9104
rect 25774 9092 25780 9104
rect 14424 9064 25780 9092
rect 14424 9052 14430 9064
rect 25774 9052 25780 9064
rect 25832 9052 25838 9104
rect 12802 8984 12808 9036
rect 12860 9024 12866 9036
rect 28534 9024 28540 9036
rect 12860 8996 28540 9024
rect 12860 8984 12866 8996
rect 28534 8984 28540 8996
rect 28592 8984 28598 9036
rect 17310 8916 17316 8968
rect 17368 8956 17374 8968
rect 30926 8956 30932 8968
rect 17368 8928 30932 8956
rect 17368 8916 17374 8928
rect 30926 8916 30932 8928
rect 30984 8916 30990 8968
rect 11238 8848 11244 8900
rect 11296 8888 11302 8900
rect 28258 8888 28264 8900
rect 11296 8860 28264 8888
rect 11296 8848 11302 8860
rect 28258 8848 28264 8860
rect 28316 8848 28322 8900
rect 8018 8780 8024 8832
rect 8076 8820 8082 8832
rect 14826 8820 14832 8832
rect 8076 8792 14832 8820
rect 8076 8780 8082 8792
rect 14826 8780 14832 8792
rect 14884 8780 14890 8832
rect 20622 8780 20628 8832
rect 20680 8820 20686 8832
rect 27430 8820 27436 8832
rect 20680 8792 27436 8820
rect 20680 8780 20686 8792
rect 27430 8780 27436 8792
rect 27488 8780 27494 8832
rect 1104 8730 33324 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 9010 8730
rect 9062 8678 9074 8730
rect 9126 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 15010 8730
rect 15062 8678 15074 8730
rect 15126 8678 15138 8730
rect 15190 8678 15202 8730
rect 15254 8678 15266 8730
rect 15318 8678 21010 8730
rect 21062 8678 21074 8730
rect 21126 8678 21138 8730
rect 21190 8678 21202 8730
rect 21254 8678 21266 8730
rect 21318 8678 27010 8730
rect 27062 8678 27074 8730
rect 27126 8678 27138 8730
rect 27190 8678 27202 8730
rect 27254 8678 27266 8730
rect 27318 8678 33010 8730
rect 33062 8678 33074 8730
rect 33126 8678 33138 8730
rect 33190 8678 33202 8730
rect 33254 8678 33266 8730
rect 33318 8678 33324 8730
rect 1104 8656 33324 8678
rect 1486 8576 1492 8628
rect 1544 8616 1550 8628
rect 1581 8619 1639 8625
rect 1581 8616 1593 8619
rect 1544 8588 1593 8616
rect 1544 8576 1550 8588
rect 1581 8585 1593 8588
rect 1627 8585 1639 8619
rect 1581 8579 1639 8585
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 3237 8619 3295 8625
rect 3237 8616 3249 8619
rect 2924 8588 3249 8616
rect 2924 8576 2930 8588
rect 3237 8585 3249 8588
rect 3283 8585 3295 8619
rect 3237 8579 3295 8585
rect 4614 8576 4620 8628
rect 4672 8616 4678 8628
rect 4801 8619 4859 8625
rect 4801 8616 4813 8619
rect 4672 8588 4813 8616
rect 4672 8576 4678 8588
rect 4801 8585 4813 8588
rect 4847 8585 4859 8619
rect 4801 8579 4859 8585
rect 6178 8576 6184 8628
rect 6236 8616 6242 8628
rect 6457 8619 6515 8625
rect 6457 8616 6469 8619
rect 6236 8588 6469 8616
rect 6236 8576 6242 8588
rect 6457 8585 6469 8588
rect 6503 8585 6515 8619
rect 6457 8579 6515 8585
rect 7742 8576 7748 8628
rect 7800 8616 7806 8628
rect 7929 8619 7987 8625
rect 7929 8616 7941 8619
rect 7800 8588 7941 8616
rect 7800 8576 7806 8588
rect 7929 8585 7941 8588
rect 7975 8585 7987 8619
rect 7929 8579 7987 8585
rect 9398 8576 9404 8628
rect 9456 8616 9462 8628
rect 9493 8619 9551 8625
rect 9493 8616 9505 8619
rect 9456 8588 9505 8616
rect 9456 8576 9462 8588
rect 9493 8585 9505 8588
rect 9539 8585 9551 8619
rect 9493 8579 9551 8585
rect 12434 8576 12440 8628
rect 12492 8616 12498 8628
rect 12621 8619 12679 8625
rect 12621 8616 12633 8619
rect 12492 8588 12633 8616
rect 12492 8576 12498 8588
rect 12621 8585 12633 8588
rect 12667 8585 12679 8619
rect 12621 8579 12679 8585
rect 13998 8576 14004 8628
rect 14056 8616 14062 8628
rect 14185 8619 14243 8625
rect 14185 8616 14197 8619
rect 14056 8588 14197 8616
rect 14056 8576 14062 8588
rect 14185 8585 14197 8588
rect 14231 8585 14243 8619
rect 14185 8579 14243 8585
rect 15562 8576 15568 8628
rect 15620 8616 15626 8628
rect 15749 8619 15807 8625
rect 15749 8616 15761 8619
rect 15620 8588 15761 8616
rect 15620 8576 15626 8588
rect 15749 8585 15761 8588
rect 15795 8585 15807 8619
rect 15749 8579 15807 8585
rect 17126 8576 17132 8628
rect 17184 8616 17190 8628
rect 17313 8619 17371 8625
rect 17313 8616 17325 8619
rect 17184 8588 17325 8616
rect 17184 8576 17190 8588
rect 17313 8585 17325 8588
rect 17359 8585 17371 8619
rect 17313 8579 17371 8585
rect 18690 8576 18696 8628
rect 18748 8616 18754 8628
rect 18877 8619 18935 8625
rect 18877 8616 18889 8619
rect 18748 8588 18889 8616
rect 18748 8576 18754 8588
rect 18877 8585 18889 8588
rect 18923 8585 18935 8619
rect 19702 8616 19708 8628
rect 18877 8579 18935 8585
rect 18984 8588 19708 8616
rect 11054 8548 11060 8560
rect 1780 8520 11060 8548
rect 1780 8489 1808 8520
rect 11054 8508 11060 8520
rect 11112 8508 11118 8560
rect 18984 8548 19012 8588
rect 19702 8576 19708 8588
rect 19760 8576 19766 8628
rect 20254 8576 20260 8628
rect 20312 8616 20318 8628
rect 20441 8619 20499 8625
rect 20441 8616 20453 8619
rect 20312 8588 20453 8616
rect 20312 8576 20318 8588
rect 20441 8585 20453 8588
rect 20487 8585 20499 8619
rect 20441 8579 20499 8585
rect 21818 8576 21824 8628
rect 21876 8616 21882 8628
rect 22005 8619 22063 8625
rect 22005 8616 22017 8619
rect 21876 8588 22017 8616
rect 21876 8576 21882 8588
rect 22005 8585 22017 8588
rect 22051 8585 22063 8619
rect 22005 8579 22063 8585
rect 23382 8576 23388 8628
rect 23440 8616 23446 8628
rect 23569 8619 23627 8625
rect 23569 8616 23581 8619
rect 23440 8588 23581 8616
rect 23440 8576 23446 8588
rect 23569 8585 23581 8588
rect 23615 8585 23627 8619
rect 23569 8579 23627 8585
rect 24946 8576 24952 8628
rect 25004 8616 25010 8628
rect 25225 8619 25283 8625
rect 25225 8616 25237 8619
rect 25004 8588 25237 8616
rect 25004 8576 25010 8588
rect 25225 8585 25237 8588
rect 25271 8585 25283 8619
rect 25225 8579 25283 8585
rect 26510 8576 26516 8628
rect 26568 8616 26574 8628
rect 27065 8619 27123 8625
rect 27065 8616 27077 8619
rect 26568 8588 27077 8616
rect 26568 8576 26574 8588
rect 27065 8585 27077 8588
rect 27111 8585 27123 8619
rect 27065 8579 27123 8585
rect 28074 8576 28080 8628
rect 28132 8616 28138 8628
rect 28261 8619 28319 8625
rect 28261 8616 28273 8619
rect 28132 8588 28273 8616
rect 28132 8576 28138 8588
rect 28261 8585 28273 8588
rect 28307 8585 28319 8619
rect 28261 8579 28319 8585
rect 29638 8576 29644 8628
rect 29696 8616 29702 8628
rect 29917 8619 29975 8625
rect 29917 8616 29929 8619
rect 29696 8588 29929 8616
rect 29696 8576 29702 8588
rect 29917 8585 29929 8588
rect 29963 8585 29975 8619
rect 29917 8579 29975 8585
rect 31110 8576 31116 8628
rect 31168 8576 31174 8628
rect 31202 8576 31208 8628
rect 31260 8616 31266 8628
rect 31481 8619 31539 8625
rect 31481 8616 31493 8619
rect 31260 8588 31493 8616
rect 31260 8576 31266 8588
rect 31481 8585 31493 8588
rect 31527 8585 31539 8619
rect 31481 8579 31539 8585
rect 32766 8576 32772 8628
rect 32824 8616 32830 8628
rect 32861 8619 32919 8625
rect 32861 8616 32873 8619
rect 32824 8588 32873 8616
rect 32824 8576 32830 8588
rect 32861 8585 32873 8588
rect 32907 8585 32919 8619
rect 32861 8579 32919 8585
rect 25314 8548 25320 8560
rect 17512 8520 19012 8548
rect 19076 8520 25320 8548
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8449 1823 8483
rect 1765 8443 1823 8449
rect 3421 8483 3479 8489
rect 3421 8449 3433 8483
rect 3467 8480 3479 8483
rect 4985 8483 5043 8489
rect 3467 8452 4936 8480
rect 3467 8449 3479 8452
rect 3421 8443 3479 8449
rect 4908 8276 4936 8452
rect 4985 8449 4997 8483
rect 5031 8449 5043 8483
rect 4985 8443 5043 8449
rect 6641 8483 6699 8489
rect 6641 8449 6653 8483
rect 6687 8480 6699 8483
rect 8018 8480 8024 8492
rect 6687 8452 8024 8480
rect 6687 8449 6699 8452
rect 6641 8443 6699 8449
rect 5000 8344 5028 8443
rect 8018 8440 8024 8452
rect 8076 8440 8082 8492
rect 8113 8483 8171 8489
rect 8113 8449 8125 8483
rect 8159 8449 8171 8483
rect 8113 8443 8171 8449
rect 9677 8483 9735 8489
rect 9677 8449 9689 8483
rect 9723 8449 9735 8483
rect 9677 8443 9735 8449
rect 8128 8344 8156 8443
rect 9692 8412 9720 8443
rect 11238 8440 11244 8492
rect 11296 8440 11302 8492
rect 12802 8440 12808 8492
rect 12860 8440 12866 8492
rect 14366 8440 14372 8492
rect 14424 8440 14430 8492
rect 15933 8483 15991 8489
rect 15933 8449 15945 8483
rect 15979 8480 15991 8483
rect 17402 8480 17408 8492
rect 15979 8452 17408 8480
rect 15979 8449 15991 8452
rect 15933 8443 15991 8449
rect 17402 8440 17408 8452
rect 17460 8440 17466 8492
rect 17512 8489 17540 8520
rect 19076 8489 19104 8520
rect 25314 8508 25320 8520
rect 25372 8508 25378 8560
rect 30650 8508 30656 8560
rect 30708 8548 30714 8560
rect 30708 8520 31708 8548
rect 30708 8508 30714 8520
rect 17497 8483 17555 8489
rect 17497 8449 17509 8483
rect 17543 8449 17555 8483
rect 17497 8443 17555 8449
rect 19061 8483 19119 8489
rect 19061 8449 19073 8483
rect 19107 8449 19119 8483
rect 19061 8443 19119 8449
rect 20622 8440 20628 8492
rect 20680 8440 20686 8492
rect 22189 8483 22247 8489
rect 22189 8449 22201 8483
rect 22235 8449 22247 8483
rect 22189 8443 22247 8449
rect 23753 8483 23811 8489
rect 23753 8449 23765 8483
rect 23799 8480 23811 8483
rect 23799 8452 24808 8480
rect 23799 8449 23811 8452
rect 23753 8443 23811 8449
rect 22204 8412 22232 8443
rect 24780 8412 24808 8452
rect 24854 8440 24860 8492
rect 24912 8480 24918 8492
rect 25041 8483 25099 8489
rect 25041 8480 25053 8483
rect 24912 8452 25053 8480
rect 24912 8440 24918 8452
rect 25041 8449 25053 8452
rect 25087 8449 25099 8483
rect 25041 8443 25099 8449
rect 27249 8483 27307 8489
rect 27249 8449 27261 8483
rect 27295 8480 27307 8483
rect 27982 8480 27988 8492
rect 27295 8452 27988 8480
rect 27295 8449 27307 8452
rect 27249 8443 27307 8449
rect 27982 8440 27988 8452
rect 28040 8440 28046 8492
rect 28445 8483 28503 8489
rect 28445 8449 28457 8483
rect 28491 8480 28503 8483
rect 28718 8480 28724 8492
rect 28491 8452 28724 8480
rect 28491 8449 28503 8452
rect 28445 8443 28503 8449
rect 28718 8440 28724 8452
rect 28776 8440 28782 8492
rect 29730 8440 29736 8492
rect 29788 8440 29794 8492
rect 30926 8440 30932 8492
rect 30984 8440 30990 8492
rect 31294 8440 31300 8492
rect 31352 8440 31358 8492
rect 31680 8489 31708 8520
rect 31665 8483 31723 8489
rect 31665 8449 31677 8483
rect 31711 8449 31723 8483
rect 31665 8443 31723 8449
rect 32309 8483 32367 8489
rect 32309 8449 32321 8483
rect 32355 8449 32367 8483
rect 32309 8443 32367 8449
rect 30834 8412 30840 8424
rect 9692 8384 22094 8412
rect 22204 8384 23789 8412
rect 24780 8384 30840 8412
rect 5000 8316 8064 8344
rect 8128 8316 10824 8344
rect 5534 8276 5540 8288
rect 4908 8248 5540 8276
rect 5534 8236 5540 8248
rect 5592 8236 5598 8288
rect 8036 8276 8064 8316
rect 9490 8276 9496 8288
rect 8036 8248 9496 8276
rect 9490 8236 9496 8248
rect 9548 8236 9554 8288
rect 10796 8276 10824 8316
rect 10870 8304 10876 8356
rect 10928 8344 10934 8356
rect 11057 8347 11115 8353
rect 11057 8344 11069 8347
rect 10928 8316 11069 8344
rect 10928 8304 10934 8316
rect 11057 8313 11069 8316
rect 11103 8313 11115 8347
rect 13814 8344 13820 8356
rect 11057 8307 11115 8313
rect 11164 8316 13820 8344
rect 11164 8276 11192 8316
rect 13814 8304 13820 8316
rect 13872 8304 13878 8356
rect 17402 8304 17408 8356
rect 17460 8344 17466 8356
rect 19426 8344 19432 8356
rect 17460 8316 19432 8344
rect 17460 8304 17466 8316
rect 19426 8304 19432 8316
rect 19484 8304 19490 8356
rect 22066 8344 22094 8384
rect 23761 8344 23789 8384
rect 30834 8372 30840 8384
rect 30892 8372 30898 8424
rect 31018 8372 31024 8424
rect 31076 8412 31082 8424
rect 32324 8412 32352 8443
rect 32398 8440 32404 8492
rect 32456 8480 32462 8492
rect 32677 8483 32735 8489
rect 32677 8480 32689 8483
rect 32456 8452 32689 8480
rect 32456 8440 32462 8452
rect 32677 8449 32689 8452
rect 32723 8449 32735 8483
rect 32677 8443 32735 8449
rect 31076 8384 32352 8412
rect 31076 8372 31082 8384
rect 29454 8344 29460 8356
rect 22066 8316 23612 8344
rect 23761 8316 29460 8344
rect 10796 8248 11192 8276
rect 23584 8276 23612 8316
rect 29454 8304 29460 8316
rect 29512 8304 29518 8356
rect 31849 8347 31907 8353
rect 31849 8313 31861 8347
rect 31895 8344 31907 8347
rect 33042 8344 33048 8356
rect 31895 8316 33048 8344
rect 31895 8313 31907 8316
rect 31849 8307 31907 8313
rect 33042 8304 33048 8316
rect 33100 8304 33106 8356
rect 24762 8276 24768 8288
rect 23584 8248 24768 8276
rect 24762 8236 24768 8248
rect 24820 8236 24826 8288
rect 32490 8236 32496 8288
rect 32548 8236 32554 8288
rect 1104 8186 33304 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 13950 8186
rect 14002 8134 14014 8186
rect 14066 8134 14078 8186
rect 14130 8134 14142 8186
rect 14194 8134 14206 8186
rect 14258 8134 19950 8186
rect 20002 8134 20014 8186
rect 20066 8134 20078 8186
rect 20130 8134 20142 8186
rect 20194 8134 20206 8186
rect 20258 8134 25950 8186
rect 26002 8134 26014 8186
rect 26066 8134 26078 8186
rect 26130 8134 26142 8186
rect 26194 8134 26206 8186
rect 26258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 33304 8186
rect 1104 8112 33304 8134
rect 17218 8032 17224 8084
rect 17276 8072 17282 8084
rect 24946 8072 24952 8084
rect 17276 8044 24952 8072
rect 17276 8032 17282 8044
rect 24946 8032 24952 8044
rect 25004 8032 25010 8084
rect 31386 8032 31392 8084
rect 31444 8032 31450 8084
rect 31754 8032 31760 8084
rect 31812 8032 31818 8084
rect 32125 8075 32183 8081
rect 32125 8041 32137 8075
rect 32171 8072 32183 8075
rect 32306 8072 32312 8084
rect 32171 8044 32312 8072
rect 32171 8041 32183 8044
rect 32125 8035 32183 8041
rect 32306 8032 32312 8044
rect 32364 8032 32370 8084
rect 16574 7964 16580 8016
rect 16632 8004 16638 8016
rect 16632 7976 32352 8004
rect 16632 7964 16638 7976
rect 1118 7896 1124 7948
rect 1176 7936 1182 7948
rect 24210 7936 24216 7948
rect 1176 7908 24216 7936
rect 1176 7896 1182 7908
rect 24210 7896 24216 7908
rect 24268 7896 24274 7948
rect 24578 7896 24584 7948
rect 24636 7936 24642 7948
rect 24636 7908 31616 7936
rect 24636 7896 24642 7908
rect 14366 7828 14372 7880
rect 14424 7868 14430 7880
rect 23014 7868 23020 7880
rect 14424 7840 23020 7868
rect 14424 7828 14430 7840
rect 23014 7828 23020 7840
rect 23072 7828 23078 7880
rect 31202 7828 31208 7880
rect 31260 7828 31266 7880
rect 31588 7877 31616 7908
rect 31573 7871 31631 7877
rect 31573 7837 31585 7871
rect 31619 7837 31631 7871
rect 31573 7831 31631 7837
rect 31662 7828 31668 7880
rect 31720 7868 31726 7880
rect 32324 7877 32352 7976
rect 31941 7871 31999 7877
rect 31941 7868 31953 7871
rect 31720 7840 31953 7868
rect 31720 7828 31726 7840
rect 31941 7837 31953 7840
rect 31987 7837 31999 7871
rect 31941 7831 31999 7837
rect 32309 7871 32367 7877
rect 32309 7837 32321 7871
rect 32355 7837 32367 7871
rect 32309 7831 32367 7837
rect 32677 7871 32735 7877
rect 32677 7837 32689 7871
rect 32723 7837 32735 7871
rect 32677 7831 32735 7837
rect 17586 7800 17592 7812
rect 6886 7772 17592 7800
rect 1394 7692 1400 7744
rect 1452 7732 1458 7744
rect 6886 7732 6914 7772
rect 17586 7760 17592 7772
rect 17644 7760 17650 7812
rect 19150 7760 19156 7812
rect 19208 7800 19214 7812
rect 32692 7800 32720 7831
rect 19208 7772 24164 7800
rect 19208 7760 19214 7772
rect 1452 7704 6914 7732
rect 1452 7692 1458 7704
rect 12342 7692 12348 7744
rect 12400 7732 12406 7744
rect 19334 7732 19340 7744
rect 12400 7704 19340 7732
rect 12400 7692 12406 7704
rect 19334 7692 19340 7704
rect 19392 7692 19398 7744
rect 24136 7732 24164 7772
rect 28966 7772 32720 7800
rect 28966 7732 28994 7772
rect 24136 7704 28994 7732
rect 32490 7692 32496 7744
rect 32548 7692 32554 7744
rect 32861 7735 32919 7741
rect 32861 7701 32873 7735
rect 32907 7732 32919 7735
rect 33594 7732 33600 7744
rect 32907 7704 33600 7732
rect 32907 7701 32919 7704
rect 32861 7695 32919 7701
rect 33594 7692 33600 7704
rect 33652 7692 33658 7744
rect 1104 7642 33324 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 9010 7642
rect 9062 7590 9074 7642
rect 9126 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 15010 7642
rect 15062 7590 15074 7642
rect 15126 7590 15138 7642
rect 15190 7590 15202 7642
rect 15254 7590 15266 7642
rect 15318 7590 21010 7642
rect 21062 7590 21074 7642
rect 21126 7590 21138 7642
rect 21190 7590 21202 7642
rect 21254 7590 21266 7642
rect 21318 7590 27010 7642
rect 27062 7590 27074 7642
rect 27126 7590 27138 7642
rect 27190 7590 27202 7642
rect 27254 7590 27266 7642
rect 27318 7590 33010 7642
rect 33062 7590 33074 7642
rect 33126 7590 33138 7642
rect 33190 7590 33202 7642
rect 33254 7590 33266 7642
rect 33318 7590 33324 7642
rect 1104 7568 33324 7590
rect 5534 7488 5540 7540
rect 5592 7528 5598 7540
rect 9309 7531 9367 7537
rect 9309 7528 9321 7531
rect 5592 7500 9321 7528
rect 5592 7488 5598 7500
rect 9309 7497 9321 7500
rect 9355 7497 9367 7531
rect 9309 7491 9367 7497
rect 11054 7488 11060 7540
rect 11112 7488 11118 7540
rect 13814 7488 13820 7540
rect 13872 7528 13878 7540
rect 14185 7531 14243 7537
rect 14185 7528 14197 7531
rect 13872 7500 14197 7528
rect 13872 7488 13878 7500
rect 14185 7497 14197 7500
rect 14231 7497 14243 7531
rect 14185 7491 14243 7497
rect 14826 7488 14832 7540
rect 14884 7488 14890 7540
rect 17586 7488 17592 7540
rect 17644 7488 17650 7540
rect 19981 7531 20039 7537
rect 19981 7497 19993 7531
rect 20027 7528 20039 7531
rect 24118 7528 24124 7540
rect 20027 7500 24124 7528
rect 20027 7497 20039 7500
rect 19981 7491 20039 7497
rect 24118 7488 24124 7500
rect 24176 7488 24182 7540
rect 24397 7531 24455 7537
rect 24397 7497 24409 7531
rect 24443 7528 24455 7531
rect 24443 7500 24716 7528
rect 24443 7497 24455 7500
rect 24397 7491 24455 7497
rect 24688 7460 24716 7500
rect 24762 7488 24768 7540
rect 24820 7488 24826 7540
rect 25314 7488 25320 7540
rect 25372 7488 25378 7540
rect 27430 7488 27436 7540
rect 27488 7528 27494 7540
rect 27709 7531 27767 7537
rect 27709 7528 27721 7531
rect 27488 7500 27721 7528
rect 27488 7488 27494 7500
rect 27709 7497 27721 7500
rect 27755 7497 27767 7531
rect 27709 7491 27767 7497
rect 27982 7488 27988 7540
rect 28040 7488 28046 7540
rect 28258 7488 28264 7540
rect 28316 7488 28322 7540
rect 28534 7488 28540 7540
rect 28592 7488 28598 7540
rect 29454 7488 29460 7540
rect 29512 7488 29518 7540
rect 30834 7488 30840 7540
rect 30892 7528 30898 7540
rect 30929 7531 30987 7537
rect 30929 7528 30941 7531
rect 30892 7500 30941 7528
rect 30892 7488 30898 7500
rect 30929 7497 30941 7500
rect 30975 7497 30987 7531
rect 30929 7491 30987 7497
rect 32493 7531 32551 7537
rect 32493 7497 32505 7531
rect 32539 7528 32551 7531
rect 33410 7528 33416 7540
rect 32539 7500 33416 7528
rect 32539 7497 32551 7500
rect 32493 7491 32551 7497
rect 33410 7488 33416 7500
rect 33468 7488 33474 7540
rect 26878 7460 26884 7472
rect 6886 7432 24072 7460
rect 24688 7432 26884 7460
rect 1210 7284 1216 7336
rect 1268 7324 1274 7336
rect 6886 7324 6914 7432
rect 9217 7395 9275 7401
rect 9217 7361 9229 7395
rect 9263 7392 9275 7395
rect 9493 7395 9551 7401
rect 9493 7392 9505 7395
rect 9263 7364 9505 7392
rect 9263 7361 9275 7364
rect 9217 7355 9275 7361
rect 9493 7361 9505 7364
rect 9539 7392 9551 7395
rect 9582 7392 9588 7404
rect 9539 7364 9588 7392
rect 9539 7361 9551 7364
rect 9493 7355 9551 7361
rect 9582 7352 9588 7364
rect 9640 7352 9646 7404
rect 11241 7395 11299 7401
rect 11241 7361 11253 7395
rect 11287 7361 11299 7395
rect 11241 7355 11299 7361
rect 1268 7296 6914 7324
rect 10873 7327 10931 7333
rect 1268 7284 1274 7296
rect 10873 7293 10885 7327
rect 10919 7324 10931 7327
rect 11256 7324 11284 7355
rect 12342 7352 12348 7404
rect 12400 7352 12406 7404
rect 14366 7352 14372 7404
rect 14424 7352 14430 7404
rect 14737 7395 14795 7401
rect 14737 7361 14749 7395
rect 14783 7392 14795 7395
rect 14918 7392 14924 7404
rect 14783 7364 14924 7392
rect 14783 7361 14795 7364
rect 14737 7355 14795 7361
rect 14918 7352 14924 7364
rect 14976 7392 14982 7404
rect 15013 7395 15071 7401
rect 15013 7392 15025 7395
rect 14976 7364 15025 7392
rect 14976 7352 14982 7364
rect 15013 7361 15025 7364
rect 15059 7361 15071 7395
rect 15013 7355 15071 7361
rect 17681 7395 17739 7401
rect 17681 7361 17693 7395
rect 17727 7392 17739 7395
rect 17773 7395 17831 7401
rect 17773 7392 17785 7395
rect 17727 7364 17785 7392
rect 17727 7361 17739 7364
rect 17681 7355 17739 7361
rect 17773 7361 17785 7364
rect 17819 7361 17831 7395
rect 17773 7355 17831 7361
rect 18046 7352 18052 7404
rect 18104 7352 18110 7404
rect 19794 7352 19800 7404
rect 19852 7352 19858 7404
rect 21818 7352 21824 7404
rect 21876 7352 21882 7404
rect 22373 7395 22431 7401
rect 22373 7361 22385 7395
rect 22419 7392 22431 7395
rect 22465 7395 22523 7401
rect 22465 7392 22477 7395
rect 22419 7364 22477 7392
rect 22419 7361 22431 7364
rect 22373 7355 22431 7361
rect 22465 7361 22477 7364
rect 22511 7361 22523 7395
rect 22465 7355 22523 7361
rect 23937 7395 23995 7401
rect 23937 7361 23949 7395
rect 23983 7361 23995 7395
rect 23937 7355 23995 7361
rect 17218 7324 17224 7336
rect 10919 7296 17224 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 17218 7284 17224 7296
rect 17276 7284 17282 7336
rect 23952 7324 23980 7355
rect 19306 7296 23980 7324
rect 24044 7324 24072 7432
rect 26878 7420 26884 7432
rect 26936 7420 26942 7472
rect 24210 7352 24216 7404
rect 24268 7352 24274 7404
rect 24489 7395 24547 7401
rect 24489 7361 24501 7395
rect 24535 7361 24547 7395
rect 24949 7395 25007 7401
rect 24489 7355 24547 7361
rect 24596 7364 24900 7392
rect 24504 7324 24532 7355
rect 24044 7296 24532 7324
rect 1670 7216 1676 7268
rect 1728 7256 1734 7268
rect 19306 7256 19334 7296
rect 24596 7256 24624 7364
rect 24762 7324 24768 7336
rect 24688 7296 24768 7324
rect 24688 7265 24716 7296
rect 24762 7284 24768 7296
rect 24820 7284 24826 7336
rect 1728 7228 19334 7256
rect 24044 7228 24624 7256
rect 24673 7259 24731 7265
rect 1728 7216 1734 7228
rect 9490 7148 9496 7200
rect 9548 7188 9554 7200
rect 12161 7191 12219 7197
rect 12161 7188 12173 7191
rect 9548 7160 12173 7188
rect 9548 7148 9554 7160
rect 12161 7157 12173 7160
rect 12207 7157 12219 7191
rect 12161 7151 12219 7157
rect 17954 7148 17960 7200
rect 18012 7148 18018 7200
rect 18230 7148 18236 7200
rect 18288 7148 18294 7200
rect 22002 7148 22008 7200
rect 22060 7148 22066 7200
rect 22278 7148 22284 7200
rect 22336 7148 22342 7200
rect 22649 7191 22707 7197
rect 22649 7157 22661 7191
rect 22695 7188 22707 7191
rect 24044 7188 24072 7228
rect 24673 7225 24685 7259
rect 24719 7225 24731 7259
rect 24872 7256 24900 7364
rect 24949 7361 24961 7395
rect 24995 7361 25007 7395
rect 24949 7355 25007 7361
rect 25501 7395 25559 7401
rect 25501 7361 25513 7395
rect 25547 7392 25559 7395
rect 25590 7392 25596 7404
rect 25547 7364 25596 7392
rect 25547 7361 25559 7364
rect 25501 7355 25559 7361
rect 24964 7324 24992 7355
rect 25590 7352 25596 7364
rect 25648 7352 25654 7404
rect 27614 7352 27620 7404
rect 27672 7392 27678 7404
rect 27893 7395 27951 7401
rect 27893 7392 27905 7395
rect 27672 7364 27905 7392
rect 27672 7352 27678 7364
rect 27893 7361 27905 7364
rect 27939 7361 27951 7395
rect 27893 7355 27951 7361
rect 27982 7352 27988 7404
rect 28040 7392 28046 7404
rect 28169 7395 28227 7401
rect 28169 7392 28181 7395
rect 28040 7364 28181 7392
rect 28040 7352 28046 7364
rect 28169 7361 28181 7364
rect 28215 7361 28227 7395
rect 28169 7355 28227 7361
rect 28442 7352 28448 7404
rect 28500 7352 28506 7404
rect 28721 7395 28779 7401
rect 28721 7361 28733 7395
rect 28767 7361 28779 7395
rect 28721 7355 28779 7361
rect 25682 7324 25688 7336
rect 24964 7296 25688 7324
rect 25682 7284 25688 7296
rect 25740 7284 25746 7336
rect 26786 7284 26792 7336
rect 26844 7324 26850 7336
rect 28736 7324 28764 7355
rect 29638 7352 29644 7404
rect 29696 7352 29702 7404
rect 30466 7352 30472 7404
rect 30524 7392 30530 7404
rect 31113 7395 31171 7401
rect 31113 7392 31125 7395
rect 30524 7364 31125 7392
rect 30524 7352 30530 7364
rect 31113 7361 31125 7364
rect 31159 7361 31171 7395
rect 31113 7355 31171 7361
rect 31386 7352 31392 7404
rect 31444 7392 31450 7404
rect 32309 7395 32367 7401
rect 32309 7392 32321 7395
rect 31444 7364 32321 7392
rect 31444 7352 31450 7364
rect 32309 7361 32321 7364
rect 32355 7361 32367 7395
rect 32309 7355 32367 7361
rect 32677 7395 32735 7401
rect 32677 7361 32689 7395
rect 32723 7361 32735 7395
rect 32677 7355 32735 7361
rect 26844 7296 28764 7324
rect 26844 7284 26850 7296
rect 30374 7284 30380 7336
rect 30432 7324 30438 7336
rect 32692 7324 32720 7355
rect 30432 7296 32720 7324
rect 30432 7284 30438 7296
rect 25866 7256 25872 7268
rect 24872 7228 25872 7256
rect 24673 7219 24731 7225
rect 25866 7216 25872 7228
rect 25924 7216 25930 7268
rect 22695 7160 24072 7188
rect 24121 7191 24179 7197
rect 22695 7157 22707 7160
rect 22649 7151 22707 7157
rect 24121 7157 24133 7191
rect 24167 7188 24179 7191
rect 30558 7188 30564 7200
rect 24167 7160 30564 7188
rect 24167 7157 24179 7160
rect 24121 7151 24179 7157
rect 30558 7148 30564 7160
rect 30616 7148 30622 7200
rect 32858 7148 32864 7200
rect 32916 7148 32922 7200
rect 1104 7098 33304 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 13950 7098
rect 14002 7046 14014 7098
rect 14066 7046 14078 7098
rect 14130 7046 14142 7098
rect 14194 7046 14206 7098
rect 14258 7046 19950 7098
rect 20002 7046 20014 7098
rect 20066 7046 20078 7098
rect 20130 7046 20142 7098
rect 20194 7046 20206 7098
rect 20258 7046 25950 7098
rect 26002 7046 26014 7098
rect 26066 7046 26078 7098
rect 26130 7046 26142 7098
rect 26194 7046 26206 7098
rect 26258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 33304 7098
rect 1104 7024 33304 7046
rect 842 6944 848 6996
rect 900 6984 906 6996
rect 21818 6984 21824 6996
rect 900 6956 21824 6984
rect 900 6944 906 6956
rect 21818 6944 21824 6956
rect 21876 6944 21882 6996
rect 24762 6944 24768 6996
rect 24820 6984 24826 6996
rect 31846 6984 31852 6996
rect 24820 6956 31852 6984
rect 24820 6944 24826 6956
rect 31846 6944 31852 6956
rect 31904 6944 31910 6996
rect 2682 6876 2688 6928
rect 2740 6916 2746 6928
rect 18046 6916 18052 6928
rect 2740 6888 18052 6916
rect 2740 6876 2746 6888
rect 18046 6876 18052 6888
rect 18104 6876 18110 6928
rect 21637 6919 21695 6925
rect 21637 6885 21649 6919
rect 21683 6885 21695 6919
rect 21637 6879 21695 6885
rect 1762 6808 1768 6860
rect 1820 6848 1826 6860
rect 1820 6820 12434 6848
rect 1820 6808 1826 6820
rect 1302 6740 1308 6792
rect 1360 6780 1366 6792
rect 12406 6780 12434 6820
rect 16482 6808 16488 6860
rect 16540 6848 16546 6860
rect 20717 6851 20775 6857
rect 20717 6848 20729 6851
rect 16540 6820 20729 6848
rect 16540 6808 16546 6820
rect 20717 6817 20729 6820
rect 20763 6848 20775 6851
rect 21652 6848 21680 6879
rect 24118 6876 24124 6928
rect 24176 6916 24182 6928
rect 30926 6916 30932 6928
rect 24176 6888 30932 6916
rect 24176 6876 24182 6888
rect 30926 6876 30932 6888
rect 30984 6876 30990 6928
rect 30374 6848 30380 6860
rect 20763 6820 21496 6848
rect 21652 6820 30380 6848
rect 20763 6817 20775 6820
rect 20717 6811 20775 6817
rect 21468 6789 21496 6820
rect 30374 6808 30380 6820
rect 30432 6808 30438 6860
rect 20257 6783 20315 6789
rect 20257 6780 20269 6783
rect 1360 6752 6914 6780
rect 12406 6752 20269 6780
rect 1360 6740 1366 6752
rect 6886 6712 6914 6752
rect 20257 6749 20269 6752
rect 20303 6749 20315 6783
rect 20257 6743 20315 6749
rect 21085 6783 21143 6789
rect 21085 6749 21097 6783
rect 21131 6780 21143 6783
rect 21177 6783 21235 6789
rect 21177 6780 21189 6783
rect 21131 6752 21189 6780
rect 21131 6749 21143 6752
rect 21085 6743 21143 6749
rect 21177 6749 21189 6752
rect 21223 6749 21235 6783
rect 21177 6743 21235 6749
rect 21453 6783 21511 6789
rect 21453 6749 21465 6783
rect 21499 6749 21511 6783
rect 21453 6743 21511 6749
rect 24581 6783 24639 6789
rect 24581 6749 24593 6783
rect 24627 6749 24639 6783
rect 24581 6743 24639 6749
rect 20993 6715 21051 6721
rect 20993 6712 21005 6715
rect 6886 6684 21005 6712
rect 20993 6681 21005 6684
rect 21039 6681 21051 6715
rect 24486 6712 24492 6724
rect 20993 6675 21051 6681
rect 21376 6684 24492 6712
rect 16114 6604 16120 6656
rect 16172 6644 16178 6656
rect 19794 6644 19800 6656
rect 16172 6616 19800 6644
rect 16172 6604 16178 6616
rect 19794 6604 19800 6616
rect 19852 6604 19858 6656
rect 20438 6604 20444 6656
rect 20496 6604 20502 6656
rect 21376 6653 21404 6684
rect 24486 6672 24492 6684
rect 24544 6672 24550 6724
rect 24596 6712 24624 6743
rect 24670 6740 24676 6792
rect 24728 6740 24734 6792
rect 25317 6783 25375 6789
rect 25317 6749 25329 6783
rect 25363 6780 25375 6783
rect 25406 6780 25412 6792
rect 25363 6752 25412 6780
rect 25363 6749 25375 6752
rect 25317 6743 25375 6749
rect 25406 6740 25412 6752
rect 25464 6740 25470 6792
rect 26237 6783 26295 6789
rect 26237 6749 26249 6783
rect 26283 6780 26295 6783
rect 26418 6780 26424 6792
rect 26283 6752 26424 6780
rect 26283 6749 26295 6752
rect 26237 6743 26295 6749
rect 26418 6740 26424 6752
rect 26476 6740 26482 6792
rect 28074 6740 28080 6792
rect 28132 6780 28138 6792
rect 28905 6783 28963 6789
rect 28905 6780 28917 6783
rect 28132 6752 28917 6780
rect 28132 6740 28138 6752
rect 28905 6749 28917 6752
rect 28951 6749 28963 6783
rect 28905 6743 28963 6749
rect 31754 6740 31760 6792
rect 31812 6780 31818 6792
rect 32309 6783 32367 6789
rect 32309 6780 32321 6783
rect 31812 6752 32321 6780
rect 31812 6740 31818 6752
rect 32309 6749 32321 6752
rect 32355 6749 32367 6783
rect 32677 6783 32735 6789
rect 32677 6780 32689 6783
rect 32309 6743 32367 6749
rect 32416 6752 32689 6780
rect 26602 6712 26608 6724
rect 24596 6684 26608 6712
rect 26602 6672 26608 6684
rect 26660 6672 26666 6724
rect 26694 6672 26700 6724
rect 26752 6712 26758 6724
rect 26752 6684 31754 6712
rect 26752 6672 26758 6684
rect 21361 6647 21419 6653
rect 21361 6613 21373 6647
rect 21407 6613 21419 6647
rect 21361 6607 21419 6613
rect 24394 6604 24400 6656
rect 24452 6604 24458 6656
rect 24854 6604 24860 6656
rect 24912 6604 24918 6656
rect 25130 6604 25136 6656
rect 25188 6604 25194 6656
rect 25774 6604 25780 6656
rect 25832 6644 25838 6656
rect 26053 6647 26111 6653
rect 26053 6644 26065 6647
rect 25832 6616 26065 6644
rect 25832 6604 25838 6616
rect 26053 6613 26065 6616
rect 26099 6613 26111 6647
rect 26053 6607 26111 6613
rect 28718 6604 28724 6656
rect 28776 6604 28782 6656
rect 31726 6644 31754 6684
rect 32416 6644 32444 6752
rect 32677 6749 32689 6752
rect 32723 6749 32735 6783
rect 32677 6743 32735 6749
rect 33410 6712 33416 6724
rect 32508 6684 33416 6712
rect 32508 6653 32536 6684
rect 33410 6672 33416 6684
rect 33468 6672 33474 6724
rect 31726 6616 32444 6644
rect 32493 6647 32551 6653
rect 32493 6613 32505 6647
rect 32539 6613 32551 6647
rect 32493 6607 32551 6613
rect 32858 6604 32864 6656
rect 32916 6604 32922 6656
rect 1104 6554 33324 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 9010 6554
rect 9062 6502 9074 6554
rect 9126 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 15010 6554
rect 15062 6502 15074 6554
rect 15126 6502 15138 6554
rect 15190 6502 15202 6554
rect 15254 6502 15266 6554
rect 15318 6502 21010 6554
rect 21062 6502 21074 6554
rect 21126 6502 21138 6554
rect 21190 6502 21202 6554
rect 21254 6502 21266 6554
rect 21318 6502 27010 6554
rect 27062 6502 27074 6554
rect 27126 6502 27138 6554
rect 27190 6502 27202 6554
rect 27254 6502 27266 6554
rect 27318 6502 33010 6554
rect 33062 6502 33074 6554
rect 33126 6502 33138 6554
rect 33190 6502 33202 6554
rect 33254 6502 33266 6554
rect 33318 6502 33324 6554
rect 1104 6480 33324 6502
rect 2590 6400 2596 6452
rect 2648 6440 2654 6452
rect 2648 6412 6914 6440
rect 2648 6400 2654 6412
rect 6886 6304 6914 6412
rect 15562 6400 15568 6452
rect 15620 6440 15626 6452
rect 15620 6412 18644 6440
rect 15620 6400 15626 6412
rect 15102 6332 15108 6384
rect 15160 6372 15166 6384
rect 18509 6375 18567 6381
rect 18509 6372 18521 6375
rect 15160 6344 18521 6372
rect 15160 6332 15166 6344
rect 18509 6341 18521 6344
rect 18555 6341 18567 6375
rect 18616 6372 18644 6412
rect 19150 6400 19156 6452
rect 19208 6400 19214 6452
rect 19702 6400 19708 6452
rect 19760 6440 19766 6452
rect 24394 6440 24400 6452
rect 19760 6412 24400 6440
rect 19760 6400 19766 6412
rect 24394 6400 24400 6412
rect 24452 6400 24458 6452
rect 24486 6400 24492 6452
rect 24544 6440 24550 6452
rect 24544 6412 25268 6440
rect 24544 6400 24550 6412
rect 18616 6344 19196 6372
rect 18509 6335 18567 6341
rect 18141 6307 18199 6313
rect 18141 6304 18153 6307
rect 6886 6276 18153 6304
rect 18141 6273 18153 6276
rect 18187 6273 18199 6307
rect 18141 6267 18199 6273
rect 18693 6307 18751 6313
rect 18693 6273 18705 6307
rect 18739 6273 18751 6307
rect 18693 6267 18751 6273
rect 2774 6196 2780 6248
rect 2832 6236 2838 6248
rect 16114 6236 16120 6248
rect 2832 6208 16120 6236
rect 2832 6196 2838 6208
rect 16114 6196 16120 6208
rect 16172 6196 16178 6248
rect 18601 6171 18659 6177
rect 18601 6137 18613 6171
rect 18647 6168 18659 6171
rect 18708 6168 18736 6267
rect 18966 6264 18972 6316
rect 19024 6264 19030 6316
rect 19168 6304 19196 6344
rect 19426 6332 19432 6384
rect 19484 6372 19490 6384
rect 25130 6372 25136 6384
rect 19484 6344 25136 6372
rect 19484 6332 19490 6344
rect 25130 6332 25136 6344
rect 25188 6332 25194 6384
rect 25240 6372 25268 6412
rect 29730 6400 29736 6452
rect 29788 6400 29794 6452
rect 32858 6400 32864 6452
rect 32916 6400 32922 6452
rect 31202 6372 31208 6384
rect 25240 6344 31208 6372
rect 31202 6332 31208 6344
rect 31260 6332 31266 6384
rect 24578 6304 24584 6316
rect 19168 6276 24584 6304
rect 24578 6264 24584 6276
rect 24636 6264 24642 6316
rect 29914 6264 29920 6316
rect 29972 6264 29978 6316
rect 32306 6264 32312 6316
rect 32364 6264 32370 6316
rect 32677 6307 32735 6313
rect 32677 6273 32689 6307
rect 32723 6273 32735 6307
rect 32677 6267 32735 6273
rect 31018 6236 31024 6248
rect 18647 6140 18736 6168
rect 18800 6208 31024 6236
rect 18647 6137 18659 6140
rect 18601 6131 18659 6137
rect 18325 6103 18383 6109
rect 18325 6069 18337 6103
rect 18371 6100 18383 6103
rect 18800 6100 18828 6208
rect 31018 6196 31024 6208
rect 31076 6196 31082 6248
rect 18877 6171 18935 6177
rect 18877 6137 18889 6171
rect 18923 6168 18935 6171
rect 32692 6168 32720 6267
rect 18923 6140 32720 6168
rect 18923 6137 18935 6140
rect 18877 6131 18935 6137
rect 18371 6072 18828 6100
rect 18371 6069 18383 6072
rect 18325 6063 18383 6069
rect 18966 6060 18972 6112
rect 19024 6100 19030 6112
rect 19245 6103 19303 6109
rect 19245 6100 19257 6103
rect 19024 6072 19257 6100
rect 19024 6060 19030 6072
rect 19245 6069 19257 6072
rect 19291 6069 19303 6103
rect 19245 6063 19303 6069
rect 32490 6060 32496 6112
rect 32548 6060 32554 6112
rect 1104 6010 33304 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 13950 6010
rect 14002 5958 14014 6010
rect 14066 5958 14078 6010
rect 14130 5958 14142 6010
rect 14194 5958 14206 6010
rect 14258 5958 19950 6010
rect 20002 5958 20014 6010
rect 20066 5958 20078 6010
rect 20130 5958 20142 6010
rect 20194 5958 20206 6010
rect 20258 5958 25950 6010
rect 26002 5958 26014 6010
rect 26066 5958 26078 6010
rect 26130 5958 26142 6010
rect 26194 5958 26206 6010
rect 26258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 33304 6010
rect 1104 5936 33304 5958
rect 17034 5856 17040 5908
rect 17092 5856 17098 5908
rect 20438 5856 20444 5908
rect 20496 5896 20502 5908
rect 30650 5896 30656 5908
rect 20496 5868 30656 5896
rect 20496 5856 20502 5868
rect 30650 5856 30656 5868
rect 30708 5856 30714 5908
rect 31021 5899 31079 5905
rect 31021 5865 31033 5899
rect 31067 5896 31079 5899
rect 31294 5896 31300 5908
rect 31067 5868 31300 5896
rect 31067 5865 31079 5868
rect 31021 5859 31079 5865
rect 31294 5856 31300 5868
rect 31352 5856 31358 5908
rect 9582 5788 9588 5840
rect 9640 5828 9646 5840
rect 24854 5828 24860 5840
rect 9640 5800 24860 5828
rect 9640 5788 9646 5800
rect 24854 5788 24860 5800
rect 24912 5788 24918 5840
rect 32858 5788 32864 5840
rect 32916 5788 32922 5840
rect 17773 5763 17831 5769
rect 17773 5760 17785 5763
rect 17512 5732 17785 5760
rect 17512 5704 17540 5732
rect 17773 5729 17785 5732
rect 17819 5729 17831 5763
rect 17773 5723 17831 5729
rect 25866 5720 25872 5772
rect 25924 5760 25930 5772
rect 25924 5732 32720 5760
rect 25924 5720 25930 5732
rect 17129 5695 17187 5701
rect 17129 5661 17141 5695
rect 17175 5692 17187 5695
rect 17221 5695 17279 5701
rect 17221 5692 17233 5695
rect 17175 5664 17233 5692
rect 17175 5661 17187 5664
rect 17129 5655 17187 5661
rect 17221 5661 17233 5664
rect 17267 5661 17279 5695
rect 17221 5655 17279 5661
rect 17494 5652 17500 5704
rect 17552 5652 17558 5704
rect 17604 5664 22094 5692
rect 17405 5559 17463 5565
rect 17405 5525 17417 5559
rect 17451 5556 17463 5559
rect 17604 5556 17632 5664
rect 22066 5624 22094 5664
rect 30834 5652 30840 5704
rect 30892 5652 30898 5704
rect 30926 5652 30932 5704
rect 30984 5692 30990 5704
rect 32692 5701 32720 5732
rect 32309 5695 32367 5701
rect 32309 5692 32321 5695
rect 30984 5664 32321 5692
rect 30984 5652 30990 5664
rect 32309 5661 32321 5664
rect 32355 5661 32367 5695
rect 32309 5655 32367 5661
rect 32677 5695 32735 5701
rect 32677 5661 32689 5695
rect 32723 5661 32735 5695
rect 32677 5655 32735 5661
rect 31662 5624 31668 5636
rect 17696 5596 19932 5624
rect 22066 5596 31668 5624
rect 17696 5565 17724 5596
rect 17451 5528 17632 5556
rect 17681 5559 17739 5565
rect 17451 5525 17463 5528
rect 17405 5519 17463 5525
rect 17681 5525 17693 5559
rect 17727 5525 17739 5559
rect 19904 5556 19932 5596
rect 31662 5584 31668 5596
rect 31720 5584 31726 5636
rect 31386 5556 31392 5568
rect 19904 5528 31392 5556
rect 17681 5519 17739 5525
rect 31386 5516 31392 5528
rect 31444 5516 31450 5568
rect 32493 5559 32551 5565
rect 32493 5525 32505 5559
rect 32539 5556 32551 5559
rect 33410 5556 33416 5568
rect 32539 5528 33416 5556
rect 32539 5525 32551 5528
rect 32493 5519 32551 5525
rect 33410 5516 33416 5528
rect 33468 5516 33474 5568
rect 1104 5466 33324 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 9010 5466
rect 9062 5414 9074 5466
rect 9126 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 15010 5466
rect 15062 5414 15074 5466
rect 15126 5414 15138 5466
rect 15190 5414 15202 5466
rect 15254 5414 15266 5466
rect 15318 5414 21010 5466
rect 21062 5414 21074 5466
rect 21126 5414 21138 5466
rect 21190 5414 21202 5466
rect 21254 5414 21266 5466
rect 21318 5414 27010 5466
rect 27062 5414 27074 5466
rect 27126 5414 27138 5466
rect 27190 5414 27202 5466
rect 27254 5414 27266 5466
rect 27318 5414 33010 5466
rect 33062 5414 33074 5466
rect 33126 5414 33138 5466
rect 33190 5414 33202 5466
rect 33254 5414 33266 5466
rect 33318 5414 33324 5466
rect 1104 5392 33324 5414
rect 13446 5352 13452 5364
rect 6886 5324 13452 5352
rect 3418 5244 3424 5296
rect 3476 5284 3482 5296
rect 6886 5284 6914 5324
rect 13446 5312 13452 5324
rect 13504 5312 13510 5364
rect 15562 5312 15568 5364
rect 15620 5312 15626 5364
rect 16390 5312 16396 5364
rect 16448 5312 16454 5364
rect 16945 5355 17003 5361
rect 16945 5321 16957 5355
rect 16991 5352 17003 5355
rect 32306 5352 32312 5364
rect 16991 5324 32312 5352
rect 16991 5321 17003 5324
rect 16945 5315 17003 5321
rect 32306 5312 32312 5324
rect 32364 5312 32370 5364
rect 32858 5312 32864 5364
rect 32916 5312 32922 5364
rect 3476 5256 6914 5284
rect 3476 5244 3482 5256
rect 7374 5244 7380 5296
rect 7432 5284 7438 5296
rect 15194 5284 15200 5296
rect 7432 5256 15200 5284
rect 7432 5244 7438 5256
rect 15194 5244 15200 5256
rect 15252 5244 15258 5296
rect 15654 5244 15660 5296
rect 15712 5284 15718 5296
rect 19426 5284 19432 5296
rect 15712 5256 19432 5284
rect 15712 5244 15718 5256
rect 19426 5244 19432 5256
rect 19484 5244 19490 5296
rect 22066 5256 32720 5284
rect 3142 5176 3148 5228
rect 3200 5216 3206 5228
rect 3200 5188 6914 5216
rect 3200 5176 3206 5188
rect 6886 5080 6914 5188
rect 10042 5176 10048 5228
rect 10100 5216 10106 5228
rect 13630 5216 13636 5228
rect 10100 5188 13636 5216
rect 10100 5176 10106 5188
rect 13630 5176 13636 5188
rect 13688 5176 13694 5228
rect 14734 5176 14740 5228
rect 14792 5216 14798 5228
rect 15289 5219 15347 5225
rect 15289 5216 15301 5219
rect 14792 5188 15301 5216
rect 14792 5176 14798 5188
rect 15289 5185 15301 5188
rect 15335 5216 15347 5219
rect 15381 5219 15439 5225
rect 15381 5216 15393 5219
rect 15335 5188 15393 5216
rect 15335 5185 15347 5188
rect 15289 5179 15347 5185
rect 15381 5185 15393 5188
rect 15427 5185 15439 5219
rect 15381 5179 15439 5185
rect 16485 5219 16543 5225
rect 16485 5185 16497 5219
rect 16531 5216 16543 5219
rect 16761 5219 16819 5225
rect 16761 5216 16773 5219
rect 16531 5188 16773 5216
rect 16531 5185 16543 5188
rect 16485 5179 16543 5185
rect 16761 5185 16773 5188
rect 16807 5185 16819 5219
rect 16761 5179 16819 5185
rect 16942 5176 16948 5228
rect 17000 5216 17006 5228
rect 17037 5219 17095 5225
rect 17037 5216 17049 5219
rect 17000 5188 17049 5216
rect 17000 5176 17006 5188
rect 17037 5185 17049 5188
rect 17083 5216 17095 5219
rect 17313 5219 17371 5225
rect 17313 5216 17325 5219
rect 17083 5188 17325 5216
rect 17083 5185 17095 5188
rect 17037 5179 17095 5185
rect 17313 5185 17325 5188
rect 17359 5185 17371 5219
rect 17313 5179 17371 5185
rect 18230 5176 18236 5228
rect 18288 5216 18294 5228
rect 22066 5216 22094 5256
rect 18288 5188 22094 5216
rect 18288 5176 18294 5188
rect 28626 5176 28632 5228
rect 28684 5216 28690 5228
rect 32692 5225 32720 5256
rect 28721 5219 28779 5225
rect 28721 5216 28733 5219
rect 28684 5188 28733 5216
rect 28684 5176 28690 5188
rect 28721 5185 28733 5188
rect 28767 5185 28779 5219
rect 28721 5179 28779 5185
rect 32309 5219 32367 5225
rect 32309 5185 32321 5219
rect 32355 5185 32367 5219
rect 32309 5179 32367 5185
rect 32677 5219 32735 5225
rect 32677 5185 32689 5219
rect 32723 5185 32735 5219
rect 32677 5179 32735 5185
rect 13262 5108 13268 5160
rect 13320 5148 13326 5160
rect 13320 5120 17908 5148
rect 13320 5108 13326 5120
rect 15470 5080 15476 5092
rect 6886 5052 15476 5080
rect 15470 5040 15476 5052
rect 15528 5040 15534 5092
rect 17221 5083 17279 5089
rect 17221 5049 17233 5083
rect 17267 5080 17279 5083
rect 17310 5080 17316 5092
rect 17267 5052 17316 5080
rect 17267 5049 17279 5052
rect 17221 5043 17279 5049
rect 17310 5040 17316 5052
rect 17368 5040 17374 5092
rect 17880 5080 17908 5120
rect 17954 5108 17960 5160
rect 18012 5148 18018 5160
rect 32324 5148 32352 5179
rect 18012 5120 32352 5148
rect 18012 5108 18018 5120
rect 21726 5080 21732 5092
rect 17880 5052 21732 5080
rect 21726 5040 21732 5052
rect 21784 5040 21790 5092
rect 28905 5083 28963 5089
rect 28905 5049 28917 5083
rect 28951 5080 28963 5083
rect 32398 5080 32404 5092
rect 28951 5052 32404 5080
rect 28951 5049 28963 5052
rect 28905 5043 28963 5049
rect 32398 5040 32404 5052
rect 32456 5040 32462 5092
rect 12066 4972 12072 5024
rect 12124 5012 12130 5024
rect 17126 5012 17132 5024
rect 12124 4984 17132 5012
rect 12124 4972 12130 4984
rect 17126 4972 17132 4984
rect 17184 4972 17190 5024
rect 32490 4972 32496 5024
rect 32548 4972 32554 5024
rect 1104 4922 33304 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 13950 4922
rect 14002 4870 14014 4922
rect 14066 4870 14078 4922
rect 14130 4870 14142 4922
rect 14194 4870 14206 4922
rect 14258 4870 19950 4922
rect 20002 4870 20014 4922
rect 20066 4870 20078 4922
rect 20130 4870 20142 4922
rect 20194 4870 20206 4922
rect 20258 4870 25950 4922
rect 26002 4870 26014 4922
rect 26066 4870 26078 4922
rect 26130 4870 26142 4922
rect 26194 4870 26206 4922
rect 26258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 33304 4922
rect 1104 4848 33304 4870
rect 3142 4768 3148 4820
rect 3200 4768 3206 4820
rect 3418 4768 3424 4820
rect 3476 4768 3482 4820
rect 7374 4768 7380 4820
rect 7432 4768 7438 4820
rect 10962 4768 10968 4820
rect 11020 4808 11026 4820
rect 11020 4780 11928 4808
rect 11020 4768 11026 4780
rect 11698 4740 11704 4752
rect 10796 4712 11704 4740
rect 6178 4672 6184 4684
rect 2976 4644 6184 4672
rect 2976 4613 3004 4644
rect 6178 4632 6184 4644
rect 6236 4632 6242 4684
rect 2961 4607 3019 4613
rect 2961 4573 2973 4607
rect 3007 4573 3019 4607
rect 2961 4567 3019 4573
rect 3237 4607 3295 4613
rect 3237 4573 3249 4607
rect 3283 4573 3295 4607
rect 3237 4567 3295 4573
rect 3789 4607 3847 4613
rect 3789 4573 3801 4607
rect 3835 4604 3847 4607
rect 5810 4604 5816 4616
rect 3835 4576 5816 4604
rect 3835 4573 3847 4576
rect 3789 4567 3847 4573
rect 3252 4536 3280 4567
rect 5810 4564 5816 4576
rect 5868 4564 5874 4616
rect 7193 4607 7251 4613
rect 7193 4573 7205 4607
rect 7239 4604 7251 4607
rect 8846 4604 8852 4616
rect 7239 4576 8852 4604
rect 7239 4573 7251 4576
rect 7193 4567 7251 4573
rect 8846 4564 8852 4576
rect 8904 4564 8910 4616
rect 10796 4613 10824 4712
rect 11698 4700 11704 4712
rect 11756 4700 11762 4752
rect 11514 4672 11520 4684
rect 11072 4644 11520 4672
rect 11072 4613 11100 4644
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 10781 4607 10839 4613
rect 10781 4573 10793 4607
rect 10827 4573 10839 4607
rect 10781 4567 10839 4573
rect 11057 4607 11115 4613
rect 11057 4573 11069 4607
rect 11103 4573 11115 4607
rect 11057 4567 11115 4573
rect 11330 4564 11336 4616
rect 11388 4564 11394 4616
rect 11900 4613 11928 4780
rect 12066 4768 12072 4820
rect 12124 4768 12130 4820
rect 13541 4811 13599 4817
rect 13541 4777 13553 4811
rect 13587 4808 13599 4811
rect 13587 4780 15148 4808
rect 13587 4777 13599 4780
rect 13541 4771 13599 4777
rect 13262 4700 13268 4752
rect 13320 4700 13326 4752
rect 11974 4632 11980 4684
rect 12032 4672 12038 4684
rect 15120 4672 15148 4780
rect 15378 4768 15384 4820
rect 15436 4768 15442 4820
rect 15930 4768 15936 4820
rect 15988 4768 15994 4820
rect 16206 4768 16212 4820
rect 16264 4768 16270 4820
rect 22002 4768 22008 4820
rect 22060 4808 22066 4820
rect 22060 4780 32720 4808
rect 22060 4768 22066 4780
rect 15197 4743 15255 4749
rect 15197 4709 15209 4743
rect 15243 4740 15255 4743
rect 16390 4740 16396 4752
rect 15243 4712 16396 4740
rect 15243 4709 15255 4712
rect 15197 4703 15255 4709
rect 16390 4700 16396 4712
rect 16448 4700 16454 4752
rect 16577 4743 16635 4749
rect 16577 4709 16589 4743
rect 16623 4740 16635 4743
rect 16623 4712 22094 4740
rect 16623 4709 16635 4712
rect 16577 4703 16635 4709
rect 20622 4672 20628 4684
rect 12032 4644 14780 4672
rect 15120 4644 20628 4672
rect 12032 4632 12038 4644
rect 11609 4607 11667 4613
rect 11609 4573 11621 4607
rect 11655 4573 11667 4607
rect 11609 4567 11667 4573
rect 11885 4607 11943 4613
rect 11885 4573 11897 4607
rect 11931 4573 11943 4607
rect 11885 4567 11943 4573
rect 5994 4536 6000 4548
rect 3252 4508 6000 4536
rect 5994 4496 6000 4508
rect 6052 4496 6058 4548
rect 11146 4496 11152 4548
rect 11204 4536 11210 4548
rect 11624 4536 11652 4567
rect 12250 4564 12256 4616
rect 12308 4564 12314 4616
rect 12526 4564 12532 4616
rect 12584 4564 12590 4616
rect 13078 4564 13084 4616
rect 13136 4564 13142 4616
rect 13354 4564 13360 4616
rect 13412 4564 13418 4616
rect 13630 4564 13636 4616
rect 13688 4564 13694 4616
rect 14752 4613 14780 4644
rect 20622 4632 20628 4644
rect 20680 4632 20686 4684
rect 22066 4672 22094 4712
rect 23198 4700 23204 4752
rect 23256 4740 23262 4752
rect 28721 4743 28779 4749
rect 28721 4740 28733 4743
rect 23256 4712 28733 4740
rect 23256 4700 23262 4712
rect 28721 4709 28733 4712
rect 28767 4709 28779 4743
rect 28721 4703 28779 4709
rect 31754 4672 31760 4684
rect 22066 4644 31760 4672
rect 31754 4632 31760 4644
rect 31812 4632 31818 4684
rect 14737 4607 14795 4613
rect 14737 4573 14749 4607
rect 14783 4573 14795 4607
rect 15013 4607 15071 4613
rect 15013 4604 15025 4607
rect 14737 4567 14795 4573
rect 14844 4576 15025 4604
rect 11204 4508 11652 4536
rect 11204 4496 11210 4508
rect 12066 4496 12072 4548
rect 12124 4536 12130 4548
rect 14844 4536 14872 4576
rect 15013 4573 15025 4576
rect 15059 4573 15071 4607
rect 15013 4567 15071 4573
rect 15381 4607 15439 4613
rect 15381 4573 15393 4607
rect 15427 4604 15439 4607
rect 15473 4607 15531 4613
rect 15473 4604 15485 4607
rect 15427 4576 15485 4604
rect 15427 4573 15439 4576
rect 15381 4567 15439 4573
rect 15473 4573 15485 4576
rect 15519 4573 15531 4607
rect 15473 4567 15531 4573
rect 15746 4564 15752 4616
rect 15804 4604 15810 4616
rect 16025 4607 16083 4613
rect 16025 4604 16037 4607
rect 15804 4576 16037 4604
rect 15804 4564 15810 4576
rect 16025 4573 16037 4576
rect 16071 4573 16083 4607
rect 16025 4567 16083 4573
rect 16301 4607 16359 4613
rect 16301 4573 16313 4607
rect 16347 4604 16359 4607
rect 16393 4607 16451 4613
rect 16393 4604 16405 4607
rect 16347 4576 16405 4604
rect 16347 4573 16359 4576
rect 16301 4567 16359 4573
rect 16393 4573 16405 4576
rect 16439 4573 16451 4607
rect 16393 4567 16451 4573
rect 25130 4564 25136 4616
rect 25188 4604 25194 4616
rect 27798 4604 27804 4616
rect 25188 4576 27804 4604
rect 25188 4564 25194 4576
rect 27798 4564 27804 4576
rect 27856 4564 27862 4616
rect 27890 4564 27896 4616
rect 27948 4564 27954 4616
rect 28258 4564 28264 4616
rect 28316 4604 28322 4616
rect 28629 4607 28687 4613
rect 28629 4604 28641 4607
rect 28316 4576 28641 4604
rect 28316 4564 28322 4576
rect 28629 4573 28641 4576
rect 28675 4573 28687 4607
rect 28629 4567 28687 4573
rect 28905 4607 28963 4613
rect 28905 4573 28917 4607
rect 28951 4573 28963 4607
rect 28905 4567 28963 4573
rect 19242 4536 19248 4548
rect 12124 4508 14872 4536
rect 14936 4508 19248 4536
rect 12124 4496 12130 4508
rect 3973 4471 4031 4477
rect 3973 4437 3985 4471
rect 4019 4468 4031 4471
rect 10134 4468 10140 4480
rect 4019 4440 10140 4468
rect 4019 4437 4031 4440
rect 3973 4431 4031 4437
rect 10134 4428 10140 4440
rect 10192 4428 10198 4480
rect 10965 4471 11023 4477
rect 10965 4437 10977 4471
rect 11011 4468 11023 4471
rect 11054 4468 11060 4480
rect 11011 4440 11060 4468
rect 11011 4437 11023 4440
rect 10965 4431 11023 4437
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 11238 4428 11244 4480
rect 11296 4428 11302 4480
rect 11517 4471 11575 4477
rect 11517 4437 11529 4471
rect 11563 4468 11575 4471
rect 11606 4468 11612 4480
rect 11563 4440 11612 4468
rect 11563 4437 11575 4440
rect 11517 4431 11575 4437
rect 11606 4428 11612 4440
rect 11664 4428 11670 4480
rect 11790 4428 11796 4480
rect 11848 4428 11854 4480
rect 12434 4428 12440 4480
rect 12492 4428 12498 4480
rect 12710 4428 12716 4480
rect 12768 4428 12774 4480
rect 13817 4471 13875 4477
rect 13817 4437 13829 4471
rect 13863 4468 13875 4471
rect 14826 4468 14832 4480
rect 13863 4440 14832 4468
rect 13863 4437 13875 4440
rect 13817 4431 13875 4437
rect 14826 4428 14832 4440
rect 14884 4428 14890 4480
rect 14936 4477 14964 4508
rect 19242 4496 19248 4508
rect 19300 4496 19306 4548
rect 27522 4496 27528 4548
rect 27580 4536 27586 4548
rect 27985 4539 28043 4545
rect 27985 4536 27997 4539
rect 27580 4508 27997 4536
rect 27580 4496 27586 4508
rect 27985 4505 27997 4508
rect 28031 4536 28043 4539
rect 28920 4536 28948 4567
rect 31846 4564 31852 4616
rect 31904 4604 31910 4616
rect 32692 4613 32720 4780
rect 32858 4700 32864 4752
rect 32916 4700 32922 4752
rect 32309 4607 32367 4613
rect 32309 4604 32321 4607
rect 31904 4576 32321 4604
rect 31904 4564 31910 4576
rect 32309 4573 32321 4576
rect 32355 4573 32367 4607
rect 32309 4567 32367 4573
rect 32677 4607 32735 4613
rect 32677 4573 32689 4607
rect 32723 4573 32735 4607
rect 32677 4567 32735 4573
rect 28031 4508 28948 4536
rect 28031 4505 28043 4508
rect 27985 4499 28043 4505
rect 14921 4471 14979 4477
rect 14921 4437 14933 4471
rect 14967 4437 14979 4471
rect 14921 4431 14979 4437
rect 15194 4428 15200 4480
rect 15252 4468 15258 4480
rect 15562 4468 15568 4480
rect 15252 4440 15568 4468
rect 15252 4428 15258 4440
rect 15562 4428 15568 4440
rect 15620 4428 15626 4480
rect 15657 4471 15715 4477
rect 15657 4437 15669 4471
rect 15703 4468 15715 4471
rect 16482 4468 16488 4480
rect 15703 4440 16488 4468
rect 15703 4437 15715 4440
rect 15657 4431 15715 4437
rect 16482 4428 16488 4440
rect 16540 4428 16546 4480
rect 24486 4428 24492 4480
rect 24544 4468 24550 4480
rect 27709 4471 27767 4477
rect 27709 4468 27721 4471
rect 24544 4440 27721 4468
rect 24544 4428 24550 4440
rect 27709 4437 27721 4440
rect 27755 4437 27767 4471
rect 27709 4431 27767 4437
rect 27798 4428 27804 4480
rect 27856 4468 27862 4480
rect 28445 4471 28503 4477
rect 28445 4468 28457 4471
rect 27856 4440 28457 4468
rect 27856 4428 27862 4440
rect 28445 4437 28457 4440
rect 28491 4437 28503 4471
rect 28445 4431 28503 4437
rect 32493 4471 32551 4477
rect 32493 4437 32505 4471
rect 32539 4468 32551 4471
rect 33410 4468 33416 4480
rect 32539 4440 33416 4468
rect 32539 4437 32551 4440
rect 32493 4431 32551 4437
rect 33410 4428 33416 4440
rect 33468 4428 33474 4480
rect 1104 4378 33324 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 9010 4378
rect 9062 4326 9074 4378
rect 9126 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 15010 4378
rect 15062 4326 15074 4378
rect 15126 4326 15138 4378
rect 15190 4326 15202 4378
rect 15254 4326 15266 4378
rect 15318 4326 21010 4378
rect 21062 4326 21074 4378
rect 21126 4326 21138 4378
rect 21190 4326 21202 4378
rect 21254 4326 21266 4378
rect 21318 4326 27010 4378
rect 27062 4326 27074 4378
rect 27126 4326 27138 4378
rect 27190 4326 27202 4378
rect 27254 4326 27266 4378
rect 27318 4326 33010 4378
rect 33062 4326 33074 4378
rect 33126 4326 33138 4378
rect 33190 4326 33202 4378
rect 33254 4326 33266 4378
rect 33318 4326 33324 4378
rect 1104 4304 33324 4326
rect 2682 4224 2688 4276
rect 2740 4224 2746 4276
rect 3145 4267 3203 4273
rect 3145 4233 3157 4267
rect 3191 4233 3203 4267
rect 3145 4227 3203 4233
rect 1949 4131 2007 4137
rect 1949 4097 1961 4131
rect 1995 4097 2007 4131
rect 1949 4091 2007 4097
rect 2225 4131 2283 4137
rect 2225 4097 2237 4131
rect 2271 4128 2283 4131
rect 2406 4128 2412 4140
rect 2271 4100 2412 4128
rect 2271 4097 2283 4100
rect 2225 4091 2283 4097
rect 1964 4060 1992 4091
rect 2406 4088 2412 4100
rect 2464 4088 2470 4140
rect 2501 4131 2559 4137
rect 2501 4097 2513 4131
rect 2547 4128 2559 4131
rect 2590 4128 2596 4140
rect 2547 4100 2596 4128
rect 2547 4097 2559 4100
rect 2501 4091 2559 4097
rect 2590 4088 2596 4100
rect 2648 4088 2654 4140
rect 2961 4131 3019 4137
rect 2961 4097 2973 4131
rect 3007 4097 3019 4131
rect 2961 4091 3019 4097
rect 2866 4060 2872 4072
rect 1964 4032 2872 4060
rect 2866 4020 2872 4032
rect 2924 4020 2930 4072
rect 2409 3995 2467 4001
rect 2409 3961 2421 3995
rect 2455 3992 2467 3995
rect 2774 3992 2780 4004
rect 2455 3964 2780 3992
rect 2455 3961 2467 3964
rect 2409 3955 2467 3961
rect 2774 3952 2780 3964
rect 2832 3952 2838 4004
rect 2976 3992 3004 4091
rect 3160 4060 3188 4227
rect 7006 4224 7012 4276
rect 7064 4224 7070 4276
rect 10778 4224 10784 4276
rect 10836 4264 10842 4276
rect 12250 4264 12256 4276
rect 10836 4236 12256 4264
rect 10836 4224 10842 4236
rect 12250 4224 12256 4236
rect 12308 4224 12314 4276
rect 12434 4224 12440 4276
rect 12492 4264 12498 4276
rect 20438 4264 20444 4276
rect 12492 4236 20444 4264
rect 12492 4224 12498 4236
rect 20438 4224 20444 4236
rect 20496 4224 20502 4276
rect 29365 4267 29423 4273
rect 29365 4264 29377 4267
rect 27172 4236 29377 4264
rect 7024 4168 8064 4196
rect 3418 4088 3424 4140
rect 3476 4088 3482 4140
rect 3694 4088 3700 4140
rect 3752 4088 3758 4140
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4097 4307 4131
rect 4249 4091 4307 4097
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4128 4675 4131
rect 6362 4128 6368 4140
rect 4663 4100 6368 4128
rect 4663 4097 4675 4100
rect 4617 4091 4675 4097
rect 4154 4060 4160 4072
rect 3160 4032 4160 4060
rect 4154 4020 4160 4032
rect 4212 4020 4218 4072
rect 4264 4060 4292 4091
rect 6362 4088 6368 4100
rect 6420 4088 6426 4140
rect 6546 4088 6552 4140
rect 6604 4088 6610 4140
rect 6825 4131 6883 4137
rect 6825 4097 6837 4131
rect 6871 4128 6883 4131
rect 7024 4128 7052 4168
rect 6871 4100 7052 4128
rect 7101 4131 7159 4137
rect 6871 4097 6883 4100
rect 6825 4091 6883 4097
rect 7101 4097 7113 4131
rect 7147 4128 7159 4131
rect 7282 4128 7288 4140
rect 7147 4100 7288 4128
rect 7147 4097 7159 4100
rect 7101 4091 7159 4097
rect 7282 4088 7288 4100
rect 7340 4088 7346 4140
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4128 7435 4131
rect 7558 4128 7564 4140
rect 7423 4100 7564 4128
rect 7423 4097 7435 4100
rect 7377 4091 7435 4097
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 7653 4131 7711 4137
rect 7653 4097 7665 4131
rect 7699 4128 7711 4131
rect 7742 4128 7748 4140
rect 7699 4100 7748 4128
rect 7699 4097 7711 4100
rect 7653 4091 7711 4097
rect 7742 4088 7748 4100
rect 7800 4088 7806 4140
rect 7834 4088 7840 4140
rect 7892 4128 7898 4140
rect 7929 4131 7987 4137
rect 7929 4128 7941 4131
rect 7892 4100 7941 4128
rect 7892 4088 7898 4100
rect 7929 4097 7941 4100
rect 7975 4097 7987 4131
rect 8036 4128 8064 4168
rect 11238 4156 11244 4208
rect 11296 4196 11302 4208
rect 13722 4196 13728 4208
rect 11296 4168 13728 4196
rect 11296 4156 11302 4168
rect 13722 4156 13728 4168
rect 13780 4156 13786 4208
rect 14826 4156 14832 4208
rect 14884 4196 14890 4208
rect 21358 4196 21364 4208
rect 14884 4168 21364 4196
rect 14884 4156 14890 4168
rect 21358 4156 21364 4168
rect 21416 4156 21422 4208
rect 27172 4196 27200 4236
rect 29365 4233 29377 4236
rect 29411 4233 29423 4267
rect 29365 4227 29423 4233
rect 27080 4168 27200 4196
rect 27632 4168 28304 4196
rect 8570 4128 8576 4140
rect 8036 4100 8576 4128
rect 7929 4091 7987 4097
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 13814 4088 13820 4140
rect 13872 4128 13878 4140
rect 14001 4131 14059 4137
rect 14001 4128 14013 4131
rect 13872 4100 14013 4128
rect 13872 4088 13878 4100
rect 14001 4097 14013 4100
rect 14047 4097 14059 4131
rect 14001 4091 14059 4097
rect 14461 4131 14519 4137
rect 14461 4097 14473 4131
rect 14507 4097 14519 4131
rect 14461 4091 14519 4097
rect 6454 4060 6460 4072
rect 4264 4032 6460 4060
rect 6454 4020 6460 4032
rect 6512 4020 6518 4072
rect 14366 4060 14372 4072
rect 7392 4032 14372 4060
rect 4801 3995 4859 4001
rect 2976 3964 4752 3992
rect 2133 3927 2191 3933
rect 2133 3893 2145 3927
rect 2179 3924 2191 3927
rect 3510 3924 3516 3936
rect 2179 3896 3516 3924
rect 2179 3893 2191 3896
rect 2133 3887 2191 3893
rect 3510 3884 3516 3896
rect 3568 3884 3574 3936
rect 3602 3884 3608 3936
rect 3660 3884 3666 3936
rect 3878 3884 3884 3936
rect 3936 3884 3942 3936
rect 4430 3884 4436 3936
rect 4488 3884 4494 3936
rect 4724 3924 4752 3964
rect 4801 3961 4813 3995
rect 4847 3992 4859 3995
rect 7392 3992 7420 4032
rect 14366 4020 14372 4032
rect 14424 4020 14430 4072
rect 4847 3964 7420 3992
rect 4847 3961 4859 3964
rect 4801 3955 4859 3961
rect 9674 3952 9680 4004
rect 9732 3992 9738 4004
rect 14476 3992 14504 4091
rect 14550 4088 14556 4140
rect 14608 4128 14614 4140
rect 15105 4131 15163 4137
rect 15105 4128 15117 4131
rect 14608 4100 15117 4128
rect 14608 4088 14614 4100
rect 15105 4097 15117 4100
rect 15151 4097 15163 4131
rect 15105 4091 15163 4097
rect 15381 4131 15439 4137
rect 15381 4097 15393 4131
rect 15427 4128 15439 4131
rect 15838 4128 15844 4140
rect 15427 4100 15844 4128
rect 15427 4097 15439 4100
rect 15381 4091 15439 4097
rect 15838 4088 15844 4100
rect 15896 4088 15902 4140
rect 22830 4088 22836 4140
rect 22888 4128 22894 4140
rect 27080 4128 27108 4168
rect 22888 4100 27108 4128
rect 27157 4131 27215 4137
rect 22888 4088 22894 4100
rect 27157 4097 27169 4131
rect 27203 4128 27215 4131
rect 27338 4128 27344 4140
rect 27203 4100 27344 4128
rect 27203 4097 27215 4100
rect 27157 4091 27215 4097
rect 27338 4088 27344 4100
rect 27396 4088 27402 4140
rect 27525 4131 27583 4137
rect 27525 4097 27537 4131
rect 27571 4128 27583 4131
rect 27632 4128 27660 4168
rect 28276 4137 28304 4168
rect 27571 4100 27660 4128
rect 27709 4131 27767 4137
rect 27571 4097 27583 4100
rect 27525 4091 27583 4097
rect 27709 4097 27721 4131
rect 27755 4128 27767 4131
rect 27985 4131 28043 4137
rect 27985 4128 27997 4131
rect 27755 4100 27997 4128
rect 27755 4097 27767 4100
rect 27709 4091 27767 4097
rect 27985 4097 27997 4100
rect 28031 4128 28043 4131
rect 28261 4131 28319 4137
rect 28031 4100 28212 4128
rect 28031 4097 28043 4100
rect 27985 4091 28043 4097
rect 21818 4060 21824 4072
rect 9732 3964 14504 3992
rect 14568 4032 21824 4060
rect 9732 3952 9738 3964
rect 5626 3924 5632 3936
rect 4724 3896 5632 3924
rect 5626 3884 5632 3896
rect 5684 3884 5690 3936
rect 6733 3927 6791 3933
rect 6733 3893 6745 3927
rect 6779 3924 6791 3927
rect 7190 3924 7196 3936
rect 6779 3896 7196 3924
rect 6779 3893 6791 3896
rect 6733 3887 6791 3893
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 7285 3927 7343 3933
rect 7285 3893 7297 3927
rect 7331 3924 7343 3927
rect 7466 3924 7472 3936
rect 7331 3896 7472 3924
rect 7331 3893 7343 3896
rect 7285 3887 7343 3893
rect 7466 3884 7472 3896
rect 7524 3884 7530 3936
rect 7561 3927 7619 3933
rect 7561 3893 7573 3927
rect 7607 3924 7619 3927
rect 7650 3924 7656 3936
rect 7607 3896 7656 3924
rect 7607 3893 7619 3896
rect 7561 3887 7619 3893
rect 7650 3884 7656 3896
rect 7708 3884 7714 3936
rect 7837 3927 7895 3933
rect 7837 3893 7849 3927
rect 7883 3924 7895 3927
rect 8018 3924 8024 3936
rect 7883 3896 8024 3924
rect 7883 3893 7895 3896
rect 7837 3887 7895 3893
rect 8018 3884 8024 3896
rect 8076 3884 8082 3936
rect 8113 3927 8171 3933
rect 8113 3893 8125 3927
rect 8159 3924 8171 3927
rect 13630 3924 13636 3936
rect 8159 3896 13636 3924
rect 8159 3893 8171 3896
rect 8113 3887 8171 3893
rect 13630 3884 13636 3896
rect 13688 3884 13694 3936
rect 14185 3927 14243 3933
rect 14185 3893 14197 3927
rect 14231 3924 14243 3927
rect 14568 3924 14596 4032
rect 21818 4020 21824 4032
rect 21876 4020 21882 4072
rect 23934 4020 23940 4072
rect 23992 4060 23998 4072
rect 27890 4060 27896 4072
rect 23992 4032 27896 4060
rect 23992 4020 23998 4032
rect 27890 4020 27896 4032
rect 27948 4020 27954 4072
rect 15565 3995 15623 4001
rect 15565 3961 15577 3995
rect 15611 3992 15623 3995
rect 22278 3992 22284 4004
rect 15611 3964 22284 3992
rect 15611 3961 15623 3964
rect 15565 3955 15623 3961
rect 22278 3952 22284 3964
rect 22336 3952 22342 4004
rect 24670 3952 24676 4004
rect 24728 3992 24734 4004
rect 28077 3995 28135 4001
rect 28077 3992 28089 3995
rect 24728 3964 28089 3992
rect 24728 3952 24734 3964
rect 28077 3961 28089 3964
rect 28123 3961 28135 3995
rect 28184 3992 28212 4100
rect 28261 4097 28273 4131
rect 28307 4097 28319 4131
rect 28261 4091 28319 4097
rect 28537 4131 28595 4137
rect 28537 4097 28549 4131
rect 28583 4128 28595 4131
rect 28813 4131 28871 4137
rect 28813 4128 28825 4131
rect 28583 4100 28825 4128
rect 28583 4097 28595 4100
rect 28537 4091 28595 4097
rect 28813 4097 28825 4100
rect 28859 4097 28871 4131
rect 28813 4091 28871 4097
rect 29089 4131 29147 4137
rect 29089 4097 29101 4131
rect 29135 4128 29147 4131
rect 29181 4131 29239 4137
rect 29181 4128 29193 4131
rect 29135 4100 29193 4128
rect 29135 4097 29147 4100
rect 29089 4091 29147 4097
rect 29181 4097 29193 4100
rect 29227 4097 29239 4131
rect 29181 4091 29239 4097
rect 29546 4088 29552 4140
rect 29604 4088 29610 4140
rect 30558 4088 30564 4140
rect 30616 4128 30622 4140
rect 32309 4131 32367 4137
rect 32309 4128 32321 4131
rect 30616 4100 32321 4128
rect 30616 4088 30622 4100
rect 32309 4097 32321 4100
rect 32355 4097 32367 4131
rect 32309 4091 32367 4097
rect 32677 4131 32735 4137
rect 32677 4097 32689 4131
rect 32723 4097 32735 4131
rect 32677 4091 32735 4097
rect 28442 4020 28448 4072
rect 28500 4020 28506 4072
rect 28902 4020 28908 4072
rect 28960 4060 28966 4072
rect 32692 4060 32720 4091
rect 28960 4032 32720 4060
rect 28960 4020 28966 4032
rect 28718 3992 28724 4004
rect 28184 3964 28724 3992
rect 28077 3955 28135 3961
rect 28718 3952 28724 3964
rect 28776 3952 28782 4004
rect 32858 3952 32864 4004
rect 32916 3952 32922 4004
rect 14231 3896 14596 3924
rect 14231 3893 14243 3896
rect 14185 3887 14243 3893
rect 14642 3884 14648 3936
rect 14700 3884 14706 3936
rect 15289 3927 15347 3933
rect 15289 3893 15301 3927
rect 15335 3924 15347 3927
rect 15654 3924 15660 3936
rect 15335 3896 15660 3924
rect 15335 3893 15347 3896
rect 15289 3887 15347 3893
rect 15654 3884 15660 3896
rect 15712 3884 15718 3936
rect 25498 3884 25504 3936
rect 25556 3924 25562 3936
rect 26973 3927 27031 3933
rect 26973 3924 26985 3927
rect 25556 3896 26985 3924
rect 25556 3884 25562 3896
rect 26973 3893 26985 3896
rect 27019 3893 27031 3927
rect 26973 3887 27031 3893
rect 27522 3884 27528 3936
rect 27580 3884 27586 3936
rect 27706 3884 27712 3936
rect 27764 3924 27770 3936
rect 27801 3927 27859 3933
rect 27801 3924 27813 3927
rect 27764 3896 27813 3924
rect 27764 3884 27770 3896
rect 27801 3893 27813 3896
rect 27847 3893 27859 3927
rect 27801 3887 27859 3893
rect 27890 3884 27896 3936
rect 27948 3924 27954 3936
rect 28629 3927 28687 3933
rect 28629 3924 28641 3927
rect 27948 3896 28641 3924
rect 27948 3884 27954 3896
rect 28629 3893 28641 3896
rect 28675 3893 28687 3927
rect 28629 3887 28687 3893
rect 28810 3884 28816 3936
rect 28868 3924 28874 3936
rect 28905 3927 28963 3933
rect 28905 3924 28917 3927
rect 28868 3896 28917 3924
rect 28868 3884 28874 3896
rect 28905 3893 28917 3896
rect 28951 3893 28963 3927
rect 28905 3887 28963 3893
rect 29178 3884 29184 3936
rect 29236 3884 29242 3936
rect 32490 3884 32496 3936
rect 32548 3884 32554 3936
rect 1104 3834 33304 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 13950 3834
rect 14002 3782 14014 3834
rect 14066 3782 14078 3834
rect 14130 3782 14142 3834
rect 14194 3782 14206 3834
rect 14258 3782 19950 3834
rect 20002 3782 20014 3834
rect 20066 3782 20078 3834
rect 20130 3782 20142 3834
rect 20194 3782 20206 3834
rect 20258 3782 25950 3834
rect 26002 3782 26014 3834
rect 26066 3782 26078 3834
rect 26130 3782 26142 3834
rect 26194 3782 26206 3834
rect 26258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 33304 3834
rect 1104 3760 33304 3782
rect 3694 3680 3700 3732
rect 3752 3720 3758 3732
rect 6730 3720 6736 3732
rect 3752 3692 6736 3720
rect 3752 3680 3758 3692
rect 6730 3680 6736 3692
rect 6788 3680 6794 3732
rect 7650 3680 7656 3732
rect 7708 3720 7714 3732
rect 18966 3720 18972 3732
rect 7708 3692 18972 3720
rect 7708 3680 7714 3692
rect 18966 3680 18972 3692
rect 19024 3680 19030 3732
rect 23753 3723 23811 3729
rect 23753 3720 23765 3723
rect 19076 3692 23765 3720
rect 3418 3612 3424 3664
rect 3476 3652 3482 3664
rect 6914 3652 6920 3664
rect 3476 3624 6920 3652
rect 3476 3612 3482 3624
rect 6914 3612 6920 3624
rect 6972 3612 6978 3664
rect 7006 3612 7012 3664
rect 7064 3652 7070 3664
rect 16574 3652 16580 3664
rect 7064 3624 16580 3652
rect 7064 3612 7070 3624
rect 16574 3612 16580 3624
rect 16632 3612 16638 3664
rect 17126 3612 17132 3664
rect 17184 3652 17190 3664
rect 19076 3652 19104 3692
rect 23753 3689 23765 3692
rect 23799 3689 23811 3723
rect 23753 3683 23811 3689
rect 24118 3680 24124 3732
rect 24176 3680 24182 3732
rect 24857 3723 24915 3729
rect 24857 3689 24869 3723
rect 24903 3720 24915 3723
rect 26050 3720 26056 3732
rect 24903 3692 26056 3720
rect 24903 3689 24915 3692
rect 24857 3683 24915 3689
rect 26050 3680 26056 3692
rect 26108 3680 26114 3732
rect 26878 3680 26884 3732
rect 26936 3720 26942 3732
rect 28902 3720 28908 3732
rect 26936 3692 28908 3720
rect 26936 3680 26942 3692
rect 28902 3680 28908 3692
rect 28960 3680 28966 3732
rect 17184 3624 19104 3652
rect 19429 3655 19487 3661
rect 17184 3612 17190 3624
rect 19429 3621 19441 3655
rect 19475 3652 19487 3655
rect 20898 3652 20904 3664
rect 19475 3624 20904 3652
rect 19475 3621 19487 3624
rect 19429 3615 19487 3621
rect 20898 3612 20904 3624
rect 20956 3612 20962 3664
rect 21177 3655 21235 3661
rect 21177 3621 21189 3655
rect 21223 3621 21235 3655
rect 21177 3615 21235 3621
rect 21453 3655 21511 3661
rect 21453 3621 21465 3655
rect 21499 3652 21511 3655
rect 24762 3652 24768 3664
rect 21499 3624 24768 3652
rect 21499 3621 21511 3624
rect 21453 3615 21511 3621
rect 2866 3544 2872 3596
rect 2924 3584 2930 3596
rect 7282 3584 7288 3596
rect 2924 3556 7288 3584
rect 2924 3544 2930 3556
rect 7282 3544 7288 3556
rect 7340 3544 7346 3596
rect 7374 3544 7380 3596
rect 7432 3584 7438 3596
rect 8386 3584 8392 3596
rect 7432 3556 8392 3584
rect 7432 3544 7438 3556
rect 8386 3544 8392 3556
rect 8444 3544 8450 3596
rect 13722 3544 13728 3596
rect 13780 3584 13786 3596
rect 19702 3584 19708 3596
rect 13780 3556 19708 3584
rect 13780 3544 13786 3556
rect 19702 3544 19708 3556
rect 19760 3544 19766 3596
rect 20714 3544 20720 3596
rect 20772 3584 20778 3596
rect 21192 3584 21220 3615
rect 24762 3612 24768 3624
rect 24820 3612 24826 3664
rect 25133 3655 25191 3661
rect 25133 3621 25145 3655
rect 25179 3652 25191 3655
rect 25179 3624 30328 3652
rect 25179 3621 25191 3624
rect 25133 3615 25191 3621
rect 22370 3584 22376 3596
rect 20772 3556 21128 3584
rect 21192 3556 22376 3584
rect 20772 3544 20778 3556
rect 2317 3519 2375 3525
rect 2317 3485 2329 3519
rect 2363 3516 2375 3519
rect 7098 3516 7104 3528
rect 2363 3488 7104 3516
rect 2363 3485 2375 3488
rect 2317 3479 2375 3485
rect 7098 3476 7104 3488
rect 7156 3476 7162 3528
rect 7193 3519 7251 3525
rect 7193 3485 7205 3519
rect 7239 3516 7251 3519
rect 8754 3516 8760 3528
rect 7239 3488 8760 3516
rect 7239 3485 7251 3488
rect 7193 3479 7251 3485
rect 8754 3476 8760 3488
rect 8812 3476 8818 3528
rect 13630 3476 13636 3528
rect 13688 3516 13694 3528
rect 17770 3516 17776 3528
rect 13688 3488 17776 3516
rect 13688 3476 13694 3488
rect 17770 3476 17776 3488
rect 17828 3476 17834 3528
rect 17865 3519 17923 3525
rect 17865 3485 17877 3519
rect 17911 3516 17923 3519
rect 17957 3519 18015 3525
rect 17957 3516 17969 3519
rect 17911 3488 17969 3516
rect 17911 3485 17923 3488
rect 17865 3479 17923 3485
rect 17957 3485 17969 3488
rect 18003 3485 18015 3519
rect 17957 3479 18015 3485
rect 19245 3519 19303 3525
rect 19245 3485 19257 3519
rect 19291 3485 19303 3519
rect 19245 3479 19303 3485
rect 20901 3519 20959 3525
rect 20901 3485 20913 3519
rect 20947 3516 20959 3519
rect 20993 3519 21051 3525
rect 20993 3516 21005 3519
rect 20947 3488 21005 3516
rect 20947 3485 20959 3488
rect 20901 3479 20959 3485
rect 20993 3485 21005 3488
rect 21039 3485 21051 3519
rect 21100 3516 21128 3556
rect 22370 3544 22376 3556
rect 22428 3544 22434 3596
rect 23382 3544 23388 3596
rect 23440 3584 23446 3596
rect 25225 3587 25283 3593
rect 25225 3584 25237 3587
rect 23440 3556 25237 3584
rect 23440 3544 23446 3556
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 21100 3488 21281 3516
rect 20993 3479 21051 3485
rect 21269 3485 21281 3488
rect 21315 3485 21327 3519
rect 21269 3479 21327 3485
rect 21554 3519 21612 3525
rect 21554 3485 21566 3519
rect 21600 3516 21612 3519
rect 21821 3519 21879 3525
rect 21600 3488 21680 3516
rect 21600 3485 21612 3488
rect 21554 3479 21612 3485
rect 2590 3408 2596 3460
rect 2648 3448 2654 3460
rect 4890 3448 4896 3460
rect 2648 3420 4896 3448
rect 2648 3408 2654 3420
rect 4890 3408 4896 3420
rect 4948 3408 4954 3460
rect 6546 3408 6552 3460
rect 6604 3448 6610 3460
rect 9398 3448 9404 3460
rect 6604 3420 9404 3448
rect 6604 3408 6610 3420
rect 9398 3408 9404 3420
rect 9456 3408 9462 3460
rect 14366 3408 14372 3460
rect 14424 3448 14430 3460
rect 17402 3448 17408 3460
rect 14424 3420 17408 3448
rect 14424 3408 14430 3420
rect 17402 3408 17408 3420
rect 17460 3408 17466 3460
rect 17494 3408 17500 3460
rect 17552 3448 17558 3460
rect 19260 3448 19288 3479
rect 19521 3451 19579 3457
rect 19521 3448 19533 3451
rect 17552 3420 19533 3448
rect 17552 3408 17558 3420
rect 19521 3417 19533 3420
rect 19567 3417 19579 3451
rect 19521 3411 19579 3417
rect 20346 3408 20352 3460
rect 20404 3448 20410 3460
rect 20404 3420 21404 3448
rect 20404 3408 20410 3420
rect 2498 3340 2504 3392
rect 2556 3340 2562 3392
rect 7374 3340 7380 3392
rect 7432 3340 7438 3392
rect 12710 3340 12716 3392
rect 12768 3380 12774 3392
rect 17586 3380 17592 3392
rect 12768 3352 17592 3380
rect 12768 3340 12774 3352
rect 17586 3340 17592 3352
rect 17644 3340 17650 3392
rect 17678 3340 17684 3392
rect 17736 3380 17742 3392
rect 17773 3383 17831 3389
rect 17773 3380 17785 3383
rect 17736 3352 17785 3380
rect 17736 3340 17742 3352
rect 17773 3349 17785 3352
rect 17819 3349 17831 3383
rect 17773 3343 17831 3349
rect 18141 3383 18199 3389
rect 18141 3349 18153 3383
rect 18187 3380 18199 3383
rect 19150 3380 19156 3392
rect 18187 3352 19156 3380
rect 18187 3349 18199 3352
rect 18141 3343 18199 3349
rect 19150 3340 19156 3352
rect 19208 3340 19214 3392
rect 19610 3340 19616 3392
rect 19668 3380 19674 3392
rect 20809 3383 20867 3389
rect 20809 3380 20821 3383
rect 19668 3352 20821 3380
rect 19668 3340 19674 3352
rect 20809 3349 20821 3352
rect 20855 3349 20867 3383
rect 21376 3380 21404 3420
rect 21652 3392 21680 3488
rect 21821 3485 21833 3519
rect 21867 3516 21879 3519
rect 21910 3516 21916 3528
rect 21867 3488 21916 3516
rect 21867 3485 21879 3488
rect 21821 3479 21879 3485
rect 21910 3476 21916 3488
rect 21968 3516 21974 3528
rect 24688 3525 24716 3556
rect 25225 3553 25237 3556
rect 25271 3553 25283 3587
rect 25225 3547 25283 3553
rect 25314 3544 25320 3596
rect 25372 3584 25378 3596
rect 26142 3584 26148 3596
rect 25372 3556 26148 3584
rect 25372 3544 25378 3556
rect 26142 3544 26148 3556
rect 26200 3544 26206 3596
rect 26786 3584 26792 3596
rect 26344 3556 26792 3584
rect 26344 3528 26372 3556
rect 26786 3544 26792 3556
rect 26844 3544 26850 3596
rect 27798 3584 27804 3596
rect 27632 3556 27804 3584
rect 22281 3519 22339 3525
rect 22281 3516 22293 3519
rect 21968 3488 22293 3516
rect 21968 3476 21974 3488
rect 22281 3485 22293 3488
rect 22327 3485 22339 3519
rect 22281 3479 22339 3485
rect 23661 3519 23719 3525
rect 23661 3485 23673 3519
rect 23707 3516 23719 3519
rect 23937 3519 23995 3525
rect 23937 3516 23949 3519
rect 23707 3488 23949 3516
rect 23707 3485 23719 3488
rect 23661 3479 23719 3485
rect 23937 3485 23949 3488
rect 23983 3485 23995 3519
rect 23937 3479 23995 3485
rect 24397 3519 24455 3525
rect 24397 3485 24409 3519
rect 24443 3485 24455 3519
rect 24397 3479 24455 3485
rect 24673 3519 24731 3525
rect 24673 3485 24685 3519
rect 24719 3485 24731 3519
rect 24673 3479 24731 3485
rect 23845 3451 23903 3457
rect 21744 3420 23796 3448
rect 21634 3380 21640 3392
rect 21376 3352 21640 3380
rect 20809 3343 20867 3349
rect 21634 3340 21640 3352
rect 21692 3340 21698 3392
rect 21744 3389 21772 3420
rect 21729 3383 21787 3389
rect 21729 3349 21741 3383
rect 21775 3349 21787 3383
rect 21729 3343 21787 3349
rect 22005 3383 22063 3389
rect 22005 3349 22017 3383
rect 22051 3380 22063 3383
rect 22094 3380 22100 3392
rect 22051 3352 22100 3380
rect 22051 3349 22063 3352
rect 22005 3343 22063 3349
rect 22094 3340 22100 3352
rect 22152 3340 22158 3392
rect 22186 3340 22192 3392
rect 22244 3340 22250 3392
rect 23566 3340 23572 3392
rect 23624 3340 23630 3392
rect 23768 3380 23796 3420
rect 23845 3417 23857 3451
rect 23891 3448 23903 3451
rect 24412 3448 24440 3479
rect 24854 3476 24860 3528
rect 24912 3516 24918 3528
rect 24949 3519 25007 3525
rect 24949 3516 24961 3519
rect 24912 3488 24961 3516
rect 24912 3476 24918 3488
rect 24949 3485 24961 3488
rect 24995 3516 25007 3519
rect 25409 3519 25467 3525
rect 25409 3516 25421 3519
rect 24995 3488 25421 3516
rect 24995 3485 25007 3488
rect 24949 3479 25007 3485
rect 25409 3485 25421 3488
rect 25455 3485 25467 3519
rect 25409 3479 25467 3485
rect 26326 3476 26332 3528
rect 26384 3476 26390 3528
rect 26510 3476 26516 3528
rect 26568 3516 26574 3528
rect 26605 3519 26663 3525
rect 26605 3516 26617 3519
rect 26568 3488 26617 3516
rect 26568 3476 26574 3488
rect 26605 3485 26617 3488
rect 26651 3485 26663 3519
rect 26605 3479 26663 3485
rect 26878 3476 26884 3528
rect 26936 3476 26942 3528
rect 27430 3476 27436 3528
rect 27488 3476 27494 3528
rect 23891 3420 24440 3448
rect 24504 3420 24992 3448
rect 23891 3417 23903 3420
rect 23845 3411 23903 3417
rect 24504 3380 24532 3420
rect 23768 3352 24532 3380
rect 24578 3340 24584 3392
rect 24636 3340 24642 3392
rect 24964 3380 24992 3420
rect 25038 3408 25044 3460
rect 25096 3448 25102 3460
rect 25096 3420 27568 3448
rect 25096 3408 25102 3420
rect 25314 3380 25320 3392
rect 24964 3352 25320 3380
rect 25314 3340 25320 3352
rect 25372 3340 25378 3392
rect 25774 3340 25780 3392
rect 25832 3380 25838 3392
rect 26421 3383 26479 3389
rect 26421 3380 26433 3383
rect 25832 3352 26433 3380
rect 25832 3340 25838 3352
rect 26421 3349 26433 3352
rect 26467 3349 26479 3383
rect 26421 3343 26479 3349
rect 26694 3340 26700 3392
rect 26752 3340 26758 3392
rect 26786 3340 26792 3392
rect 26844 3380 26850 3392
rect 27540 3389 27568 3420
rect 27249 3383 27307 3389
rect 27249 3380 27261 3383
rect 26844 3352 27261 3380
rect 26844 3340 26850 3352
rect 27249 3349 27261 3352
rect 27295 3349 27307 3383
rect 27249 3343 27307 3349
rect 27525 3383 27583 3389
rect 27525 3349 27537 3383
rect 27571 3349 27583 3383
rect 27632 3380 27660 3556
rect 27798 3544 27804 3556
rect 27856 3544 27862 3596
rect 27709 3519 27767 3525
rect 27709 3485 27721 3519
rect 27755 3516 27767 3519
rect 27890 3516 27896 3528
rect 27755 3488 27896 3516
rect 27755 3485 27767 3488
rect 27709 3479 27767 3485
rect 27890 3476 27896 3488
rect 27948 3476 27954 3528
rect 28169 3519 28227 3525
rect 28169 3485 28181 3519
rect 28215 3516 28227 3519
rect 28350 3516 28356 3528
rect 28215 3488 28356 3516
rect 28215 3485 28227 3488
rect 28169 3479 28227 3485
rect 27801 3451 27859 3457
rect 27801 3417 27813 3451
rect 27847 3448 27859 3451
rect 28184 3448 28212 3479
rect 28350 3476 28356 3488
rect 28408 3476 28414 3528
rect 28445 3519 28503 3525
rect 28445 3485 28457 3519
rect 28491 3516 28503 3519
rect 28537 3519 28595 3525
rect 28537 3516 28549 3519
rect 28491 3488 28549 3516
rect 28491 3485 28503 3488
rect 28445 3479 28503 3485
rect 28537 3485 28549 3488
rect 28583 3485 28595 3519
rect 28537 3479 28595 3485
rect 27847 3420 28212 3448
rect 30300 3448 30328 3624
rect 32858 3612 32864 3664
rect 32916 3612 32922 3664
rect 30374 3544 30380 3596
rect 30432 3584 30438 3596
rect 30432 3556 32720 3584
rect 30432 3544 30438 3556
rect 32692 3525 32720 3556
rect 32309 3519 32367 3525
rect 32309 3485 32321 3519
rect 32355 3485 32367 3519
rect 32309 3479 32367 3485
rect 32677 3519 32735 3525
rect 32677 3485 32689 3519
rect 32723 3485 32735 3519
rect 32677 3479 32735 3485
rect 32324 3448 32352 3479
rect 30300 3420 32352 3448
rect 27847 3417 27859 3420
rect 27801 3411 27859 3417
rect 27985 3383 28043 3389
rect 27985 3380 27997 3383
rect 27632 3352 27997 3380
rect 27525 3343 27583 3349
rect 27985 3349 27997 3352
rect 28031 3349 28043 3383
rect 27985 3343 28043 3349
rect 28166 3340 28172 3392
rect 28224 3380 28230 3392
rect 28261 3383 28319 3389
rect 28261 3380 28273 3383
rect 28224 3352 28273 3380
rect 28224 3340 28230 3352
rect 28261 3349 28273 3352
rect 28307 3349 28319 3383
rect 28261 3343 28319 3349
rect 28534 3340 28540 3392
rect 28592 3340 28598 3392
rect 32493 3383 32551 3389
rect 32493 3349 32505 3383
rect 32539 3380 32551 3383
rect 33410 3380 33416 3392
rect 32539 3352 33416 3380
rect 32539 3349 32551 3352
rect 32493 3343 32551 3349
rect 33410 3340 33416 3352
rect 33468 3340 33474 3392
rect 1104 3290 33324 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 9010 3290
rect 9062 3238 9074 3290
rect 9126 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 15010 3290
rect 15062 3238 15074 3290
rect 15126 3238 15138 3290
rect 15190 3238 15202 3290
rect 15254 3238 15266 3290
rect 15318 3238 21010 3290
rect 21062 3238 21074 3290
rect 21126 3238 21138 3290
rect 21190 3238 21202 3290
rect 21254 3238 21266 3290
rect 21318 3238 27010 3290
rect 27062 3238 27074 3290
rect 27126 3238 27138 3290
rect 27190 3238 27202 3290
rect 27254 3238 27266 3290
rect 27318 3238 33010 3290
rect 33062 3238 33074 3290
rect 33126 3238 33138 3290
rect 33190 3238 33202 3290
rect 33254 3238 33266 3290
rect 33318 3238 33324 3290
rect 1104 3216 33324 3238
rect 2406 3136 2412 3188
rect 2464 3176 2470 3188
rect 4522 3176 4528 3188
rect 2464 3148 4528 3176
rect 2464 3136 2470 3148
rect 4522 3136 4528 3148
rect 4580 3136 4586 3188
rect 10134 3136 10140 3188
rect 10192 3176 10198 3188
rect 15930 3176 15936 3188
rect 10192 3148 15936 3176
rect 10192 3136 10198 3148
rect 15930 3136 15936 3148
rect 15988 3136 15994 3188
rect 17586 3136 17592 3188
rect 17644 3176 17650 3188
rect 17644 3148 20576 3176
rect 17644 3136 17650 3148
rect 11790 3068 11796 3120
rect 11848 3108 11854 3120
rect 11848 3080 20116 3108
rect 11848 3068 11854 3080
rect 15470 3000 15476 3052
rect 15528 3000 15534 3052
rect 15841 3043 15899 3049
rect 15841 3009 15853 3043
rect 15887 3009 15899 3043
rect 15841 3003 15899 3009
rect 3878 2932 3884 2984
rect 3936 2972 3942 2984
rect 15856 2972 15884 3003
rect 16022 3000 16028 3052
rect 16080 3040 16086 3052
rect 16209 3043 16267 3049
rect 16209 3040 16221 3043
rect 16080 3012 16221 3040
rect 16080 3000 16086 3012
rect 16209 3009 16221 3012
rect 16255 3009 16267 3043
rect 16209 3003 16267 3009
rect 16758 3000 16764 3052
rect 16816 3000 16822 3052
rect 17129 3043 17187 3049
rect 17129 3009 17141 3043
rect 17175 3009 17187 3043
rect 17129 3003 17187 3009
rect 15930 2972 15936 2984
rect 3936 2944 14964 2972
rect 15856 2944 15936 2972
rect 3936 2932 3942 2944
rect 2682 2864 2688 2916
rect 2740 2904 2746 2916
rect 14826 2904 14832 2916
rect 2740 2876 14832 2904
rect 2740 2864 2746 2876
rect 14826 2864 14832 2876
rect 14884 2864 14890 2916
rect 14936 2904 14964 2944
rect 15930 2932 15936 2944
rect 15988 2932 15994 2984
rect 17144 2972 17172 3003
rect 17402 3000 17408 3052
rect 17460 3040 17466 3052
rect 17497 3043 17555 3049
rect 17497 3040 17509 3043
rect 17460 3012 17509 3040
rect 17460 3000 17466 3012
rect 17497 3009 17509 3012
rect 17543 3009 17555 3043
rect 17497 3003 17555 3009
rect 18966 3000 18972 3052
rect 19024 3000 19030 3052
rect 19242 3000 19248 3052
rect 19300 3040 19306 3052
rect 19337 3043 19395 3049
rect 19337 3040 19349 3043
rect 19300 3012 19349 3040
rect 19300 3000 19306 3012
rect 19337 3009 19349 3012
rect 19383 3009 19395 3043
rect 19337 3003 19395 3009
rect 19702 3000 19708 3052
rect 19760 3000 19766 3052
rect 20088 3049 20116 3080
rect 20073 3043 20131 3049
rect 20073 3009 20085 3043
rect 20119 3009 20131 3043
rect 20073 3003 20131 3009
rect 20438 3000 20444 3052
rect 20496 3000 20502 3052
rect 20548 3040 20576 3148
rect 22002 3136 22008 3188
rect 22060 3176 22066 3188
rect 22649 3179 22707 3185
rect 22649 3176 22661 3179
rect 22060 3148 22661 3176
rect 22060 3136 22066 3148
rect 22649 3145 22661 3148
rect 22695 3145 22707 3179
rect 22649 3139 22707 3145
rect 23658 3136 23664 3188
rect 23716 3176 23722 3188
rect 24489 3179 24547 3185
rect 24489 3176 24501 3179
rect 23716 3148 24501 3176
rect 23716 3136 23722 3148
rect 24489 3145 24501 3148
rect 24535 3145 24547 3179
rect 24489 3139 24547 3145
rect 24762 3136 24768 3188
rect 24820 3176 24826 3188
rect 25593 3179 25651 3185
rect 25593 3176 25605 3179
rect 24820 3148 25605 3176
rect 24820 3136 24826 3148
rect 25593 3145 25605 3148
rect 25639 3145 25651 3179
rect 25593 3139 25651 3145
rect 27062 3136 27068 3188
rect 27120 3176 27126 3188
rect 27522 3176 27528 3188
rect 27120 3148 27528 3176
rect 27120 3136 27126 3148
rect 27522 3136 27528 3148
rect 27580 3136 27586 3188
rect 27617 3179 27675 3185
rect 27617 3145 27629 3179
rect 27663 3145 27675 3179
rect 27617 3139 27675 3145
rect 27632 3108 27660 3139
rect 27798 3136 27804 3188
rect 27856 3136 27862 3188
rect 32858 3136 32864 3188
rect 32916 3136 32922 3188
rect 27816 3108 27844 3136
rect 24320 3080 27660 3108
rect 27724 3080 27844 3108
rect 20809 3043 20867 3049
rect 20809 3040 20821 3043
rect 20548 3012 20821 3040
rect 20809 3009 20821 3012
rect 20855 3009 20867 3043
rect 20809 3003 20867 3009
rect 21177 3043 21235 3049
rect 21177 3009 21189 3043
rect 21223 3009 21235 3043
rect 21177 3003 21235 3009
rect 16040 2944 17172 2972
rect 16040 2904 16068 2944
rect 17218 2932 17224 2984
rect 17276 2972 17282 2984
rect 20346 2972 20352 2984
rect 17276 2944 20352 2972
rect 17276 2932 17282 2944
rect 20346 2932 20352 2944
rect 20404 2932 20410 2984
rect 20622 2932 20628 2984
rect 20680 2972 20686 2984
rect 21192 2972 21220 3003
rect 21818 3000 21824 3052
rect 21876 3000 21882 3052
rect 22189 3043 22247 3049
rect 22189 3009 22201 3043
rect 22235 3040 22247 3043
rect 22278 3040 22284 3052
rect 22235 3012 22284 3040
rect 22235 3009 22247 3012
rect 22189 3003 22247 3009
rect 22278 3000 22284 3012
rect 22336 3000 22342 3052
rect 22830 3000 22836 3052
rect 22888 3000 22894 3052
rect 23198 3000 23204 3052
rect 23256 3000 23262 3052
rect 23569 3043 23627 3049
rect 23569 3009 23581 3043
rect 23615 3040 23627 3043
rect 23615 3012 23888 3040
rect 23615 3009 23627 3012
rect 23569 3003 23627 3009
rect 20680 2944 21220 2972
rect 20680 2932 20686 2944
rect 22922 2932 22928 2984
rect 22980 2972 22986 2984
rect 23860 2972 23888 3012
rect 23934 3000 23940 3052
rect 23992 3000 23998 3052
rect 24320 3049 24348 3080
rect 24305 3043 24363 3049
rect 24305 3009 24317 3043
rect 24351 3009 24363 3043
rect 24305 3003 24363 3009
rect 24670 3000 24676 3052
rect 24728 3000 24734 3052
rect 25038 3000 25044 3052
rect 25096 3000 25102 3052
rect 25409 3044 25467 3049
rect 25498 3044 25504 3052
rect 25409 3043 25504 3044
rect 25409 3009 25421 3043
rect 25455 3016 25504 3043
rect 25455 3009 25467 3016
rect 25409 3003 25467 3009
rect 25498 3000 25504 3016
rect 25556 3000 25562 3052
rect 25774 3000 25780 3052
rect 25832 3000 25838 3052
rect 27724 2972 27752 3080
rect 28442 3068 28448 3120
rect 28500 3108 28506 3120
rect 28500 3080 32352 3108
rect 28500 3068 28506 3080
rect 27798 3000 27804 3052
rect 27856 3000 27862 3052
rect 31662 3000 31668 3052
rect 31720 3000 31726 3052
rect 32324 3049 32352 3080
rect 32309 3043 32367 3049
rect 32309 3009 32321 3043
rect 32355 3009 32367 3043
rect 32309 3003 32367 3009
rect 32677 3043 32735 3049
rect 32677 3009 32689 3043
rect 32723 3009 32735 3043
rect 32677 3003 32735 3009
rect 22980 2944 23796 2972
rect 23860 2944 27752 2972
rect 22980 2932 22986 2944
rect 14936 2876 16068 2904
rect 16574 2864 16580 2916
rect 16632 2904 16638 2916
rect 17770 2904 17776 2916
rect 16632 2876 17776 2904
rect 16632 2864 16638 2876
rect 17770 2864 17776 2876
rect 17828 2864 17834 2916
rect 17862 2864 17868 2916
rect 17920 2904 17926 2916
rect 19058 2904 19064 2916
rect 17920 2876 19064 2904
rect 17920 2864 17926 2876
rect 19058 2864 19064 2876
rect 19116 2864 19122 2916
rect 19334 2864 19340 2916
rect 19392 2904 19398 2916
rect 19702 2904 19708 2916
rect 19392 2876 19708 2904
rect 19392 2864 19398 2876
rect 19702 2864 19708 2876
rect 19760 2864 19766 2916
rect 19794 2864 19800 2916
rect 19852 2904 19858 2916
rect 20257 2907 20315 2913
rect 20257 2904 20269 2907
rect 19852 2876 20269 2904
rect 19852 2864 19858 2876
rect 20257 2873 20269 2876
rect 20303 2873 20315 2907
rect 20257 2867 20315 2873
rect 20530 2864 20536 2916
rect 20588 2904 20594 2916
rect 20993 2907 21051 2913
rect 20993 2904 21005 2907
rect 20588 2876 21005 2904
rect 20588 2864 20594 2876
rect 20993 2873 21005 2876
rect 21039 2873 21051 2907
rect 20993 2867 21051 2873
rect 21634 2864 21640 2916
rect 21692 2904 21698 2916
rect 22373 2907 22431 2913
rect 22373 2904 22385 2907
rect 21692 2876 22385 2904
rect 21692 2864 21698 2876
rect 22373 2873 22385 2876
rect 22419 2873 22431 2907
rect 22373 2867 22431 2873
rect 22462 2864 22468 2916
rect 22520 2904 22526 2916
rect 23017 2907 23075 2913
rect 23017 2904 23029 2907
rect 22520 2876 23029 2904
rect 22520 2864 22526 2876
rect 23017 2873 23029 2876
rect 23063 2873 23075 2907
rect 23017 2867 23075 2873
rect 23290 2864 23296 2916
rect 23348 2904 23354 2916
rect 23768 2913 23796 2944
rect 23753 2907 23811 2913
rect 23348 2876 23520 2904
rect 23348 2864 23354 2876
rect 10594 2796 10600 2848
rect 10652 2836 10658 2848
rect 12526 2836 12532 2848
rect 10652 2808 12532 2836
rect 10652 2796 10658 2808
rect 12526 2796 12532 2808
rect 12584 2796 12590 2848
rect 15378 2796 15384 2848
rect 15436 2836 15442 2848
rect 15657 2839 15715 2845
rect 15657 2836 15669 2839
rect 15436 2808 15669 2836
rect 15436 2796 15442 2808
rect 15657 2805 15669 2808
rect 15703 2805 15715 2839
rect 15657 2799 15715 2805
rect 15746 2796 15752 2848
rect 15804 2836 15810 2848
rect 16025 2839 16083 2845
rect 16025 2836 16037 2839
rect 15804 2808 16037 2836
rect 15804 2796 15810 2808
rect 16025 2805 16037 2808
rect 16071 2805 16083 2839
rect 16025 2799 16083 2805
rect 16114 2796 16120 2848
rect 16172 2836 16178 2848
rect 16393 2839 16451 2845
rect 16393 2836 16405 2839
rect 16172 2808 16405 2836
rect 16172 2796 16178 2808
rect 16393 2805 16405 2808
rect 16439 2805 16451 2839
rect 16393 2799 16451 2805
rect 16666 2796 16672 2848
rect 16724 2836 16730 2848
rect 16945 2839 17003 2845
rect 16945 2836 16957 2839
rect 16724 2808 16957 2836
rect 16724 2796 16730 2808
rect 16945 2805 16957 2808
rect 16991 2805 17003 2839
rect 16945 2799 17003 2805
rect 17034 2796 17040 2848
rect 17092 2836 17098 2848
rect 17313 2839 17371 2845
rect 17313 2836 17325 2839
rect 17092 2808 17325 2836
rect 17092 2796 17098 2808
rect 17313 2805 17325 2808
rect 17359 2805 17371 2839
rect 17313 2799 17371 2805
rect 17402 2796 17408 2848
rect 17460 2836 17466 2848
rect 17681 2839 17739 2845
rect 17681 2836 17693 2839
rect 17460 2808 17693 2836
rect 17460 2796 17466 2808
rect 17681 2805 17693 2808
rect 17727 2805 17739 2839
rect 17681 2799 17739 2805
rect 18874 2796 18880 2848
rect 18932 2836 18938 2848
rect 19153 2839 19211 2845
rect 19153 2836 19165 2839
rect 18932 2808 19165 2836
rect 18932 2796 18938 2808
rect 19153 2805 19165 2808
rect 19199 2805 19211 2839
rect 19153 2799 19211 2805
rect 19242 2796 19248 2848
rect 19300 2836 19306 2848
rect 19521 2839 19579 2845
rect 19521 2836 19533 2839
rect 19300 2808 19533 2836
rect 19300 2796 19306 2808
rect 19521 2805 19533 2808
rect 19567 2805 19579 2839
rect 19521 2799 19579 2805
rect 19610 2796 19616 2848
rect 19668 2836 19674 2848
rect 19889 2839 19947 2845
rect 19889 2836 19901 2839
rect 19668 2808 19901 2836
rect 19668 2796 19674 2808
rect 19889 2805 19901 2808
rect 19935 2805 19947 2839
rect 19889 2799 19947 2805
rect 20346 2796 20352 2848
rect 20404 2836 20410 2848
rect 20625 2839 20683 2845
rect 20625 2836 20637 2839
rect 20404 2808 20637 2836
rect 20404 2796 20410 2808
rect 20625 2805 20637 2808
rect 20671 2805 20683 2839
rect 20625 2799 20683 2805
rect 20714 2796 20720 2848
rect 20772 2836 20778 2848
rect 21361 2839 21419 2845
rect 21361 2836 21373 2839
rect 20772 2808 21373 2836
rect 20772 2796 20778 2808
rect 21361 2805 21373 2808
rect 21407 2805 21419 2839
rect 21361 2799 21419 2805
rect 21450 2796 21456 2848
rect 21508 2836 21514 2848
rect 22005 2839 22063 2845
rect 22005 2836 22017 2839
rect 21508 2808 22017 2836
rect 21508 2796 21514 2808
rect 22005 2805 22017 2808
rect 22051 2805 22063 2839
rect 22005 2799 22063 2805
rect 22738 2796 22744 2848
rect 22796 2836 22802 2848
rect 23385 2839 23443 2845
rect 23385 2836 23397 2839
rect 22796 2808 23397 2836
rect 22796 2796 22802 2808
rect 23385 2805 23397 2808
rect 23431 2805 23443 2839
rect 23492 2836 23520 2876
rect 23753 2873 23765 2907
rect 23799 2873 23811 2907
rect 23753 2867 23811 2873
rect 24026 2864 24032 2916
rect 24084 2904 24090 2916
rect 24857 2907 24915 2913
rect 24857 2904 24869 2907
rect 24084 2876 24869 2904
rect 24084 2864 24090 2876
rect 24857 2873 24869 2876
rect 24903 2873 24915 2907
rect 25225 2907 25283 2913
rect 25225 2904 25237 2907
rect 24857 2867 24915 2873
rect 24964 2876 25237 2904
rect 24121 2839 24179 2845
rect 24121 2836 24133 2839
rect 23492 2808 24133 2836
rect 23385 2799 23443 2805
rect 24121 2805 24133 2808
rect 24167 2805 24179 2839
rect 24121 2799 24179 2805
rect 24394 2796 24400 2848
rect 24452 2836 24458 2848
rect 24964 2836 24992 2876
rect 25225 2873 25237 2876
rect 25271 2873 25283 2907
rect 25225 2867 25283 2873
rect 28258 2864 28264 2916
rect 28316 2904 28322 2916
rect 32692 2904 32720 3003
rect 28316 2876 32720 2904
rect 28316 2864 28322 2876
rect 24452 2808 24992 2836
rect 24452 2796 24458 2808
rect 25774 2796 25780 2848
rect 25832 2836 25838 2848
rect 28810 2836 28816 2848
rect 25832 2808 28816 2836
rect 25832 2796 25838 2808
rect 28810 2796 28816 2808
rect 28868 2796 28874 2848
rect 31849 2839 31907 2845
rect 31849 2805 31861 2839
rect 31895 2836 31907 2839
rect 32398 2836 32404 2848
rect 31895 2808 32404 2836
rect 31895 2805 31907 2808
rect 31849 2799 31907 2805
rect 32398 2796 32404 2808
rect 32456 2796 32462 2848
rect 32490 2796 32496 2848
rect 32548 2796 32554 2848
rect 1104 2746 33304 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 13950 2746
rect 14002 2694 14014 2746
rect 14066 2694 14078 2746
rect 14130 2694 14142 2746
rect 14194 2694 14206 2746
rect 14258 2694 19950 2746
rect 20002 2694 20014 2746
rect 20066 2694 20078 2746
rect 20130 2694 20142 2746
rect 20194 2694 20206 2746
rect 20258 2694 25950 2746
rect 26002 2694 26014 2746
rect 26066 2694 26078 2746
rect 26130 2694 26142 2746
rect 26194 2694 26206 2746
rect 26258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 33304 2746
rect 1104 2672 33304 2694
rect 3602 2592 3608 2644
rect 3660 2632 3666 2644
rect 11054 2632 11060 2644
rect 3660 2604 11060 2632
rect 3660 2592 3666 2604
rect 11054 2592 11060 2604
rect 11112 2592 11118 2644
rect 15470 2632 15476 2644
rect 11164 2604 15476 2632
rect 2774 2524 2780 2576
rect 2832 2564 2838 2576
rect 11164 2564 11192 2604
rect 15470 2592 15476 2604
rect 15528 2592 15534 2644
rect 18506 2592 18512 2644
rect 18564 2632 18570 2644
rect 19429 2635 19487 2641
rect 19429 2632 19441 2635
rect 18564 2604 19441 2632
rect 18564 2592 18570 2604
rect 19429 2601 19441 2604
rect 19475 2601 19487 2635
rect 19429 2595 19487 2601
rect 20162 2592 20168 2644
rect 20220 2632 20226 2644
rect 21269 2635 21327 2641
rect 21269 2632 21281 2635
rect 20220 2604 21281 2632
rect 20220 2592 20226 2604
rect 21269 2601 21281 2604
rect 21315 2601 21327 2635
rect 21269 2595 21327 2601
rect 21818 2592 21824 2644
rect 21876 2632 21882 2644
rect 21876 2604 22140 2632
rect 21876 2592 21882 2604
rect 2832 2536 11192 2564
rect 14921 2567 14979 2573
rect 2832 2524 2838 2536
rect 14921 2533 14933 2567
rect 14967 2564 14979 2567
rect 15562 2564 15568 2576
rect 14967 2536 15568 2564
rect 14967 2533 14979 2536
rect 14921 2527 14979 2533
rect 15562 2524 15568 2536
rect 15620 2524 15626 2576
rect 16025 2567 16083 2573
rect 16025 2533 16037 2567
rect 16071 2564 16083 2567
rect 16482 2564 16488 2576
rect 16071 2536 16488 2564
rect 16071 2533 16083 2536
rect 16025 2527 16083 2533
rect 16482 2524 16488 2536
rect 16540 2524 16546 2576
rect 18138 2524 18144 2576
rect 18196 2564 18202 2576
rect 18969 2567 19027 2573
rect 18969 2564 18981 2567
rect 18196 2536 18981 2564
rect 18196 2524 18202 2536
rect 18969 2533 18981 2536
rect 19015 2533 19027 2567
rect 18969 2527 19027 2533
rect 19886 2524 19892 2576
rect 19944 2564 19950 2576
rect 20533 2567 20591 2573
rect 20533 2564 20545 2567
rect 19944 2536 20545 2564
rect 19944 2524 19950 2536
rect 20533 2533 20545 2536
rect 20579 2533 20591 2567
rect 20533 2527 20591 2533
rect 20898 2524 20904 2576
rect 20956 2564 20962 2576
rect 22005 2567 22063 2573
rect 22005 2564 22017 2567
rect 20956 2536 22017 2564
rect 20956 2524 20962 2536
rect 22005 2533 22017 2536
rect 22051 2533 22063 2567
rect 22005 2527 22063 2533
rect 3510 2456 3516 2508
rect 3568 2496 3574 2508
rect 3568 2468 15884 2496
rect 3568 2456 3574 2468
rect 10410 2388 10416 2440
rect 10468 2428 10474 2440
rect 13354 2428 13360 2440
rect 10468 2400 13360 2428
rect 10468 2388 10474 2400
rect 13354 2388 13360 2400
rect 13412 2388 13418 2440
rect 13446 2388 13452 2440
rect 13504 2428 13510 2440
rect 14737 2431 14795 2437
rect 14737 2428 14749 2431
rect 13504 2400 14749 2428
rect 13504 2388 13510 2400
rect 14737 2397 14749 2400
rect 14783 2397 14795 2431
rect 14737 2391 14795 2397
rect 15105 2431 15163 2437
rect 15105 2397 15117 2431
rect 15151 2397 15163 2431
rect 15105 2391 15163 2397
rect 4154 2320 4160 2372
rect 4212 2360 4218 2372
rect 15120 2360 15148 2391
rect 15470 2388 15476 2440
rect 15528 2388 15534 2440
rect 15856 2437 15884 2468
rect 16298 2456 16304 2508
rect 16356 2496 16362 2508
rect 16356 2468 17724 2496
rect 16356 2456 16362 2468
rect 15841 2431 15899 2437
rect 15841 2397 15853 2431
rect 15887 2397 15899 2431
rect 15841 2391 15899 2397
rect 16206 2388 16212 2440
rect 16264 2388 16270 2440
rect 16942 2388 16948 2440
rect 17000 2388 17006 2440
rect 17310 2388 17316 2440
rect 17368 2388 17374 2440
rect 17696 2437 17724 2468
rect 17770 2456 17776 2508
rect 17828 2496 17834 2508
rect 17828 2468 18828 2496
rect 17828 2456 17834 2468
rect 17681 2431 17739 2437
rect 17681 2397 17693 2431
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 18046 2388 18052 2440
rect 18104 2388 18110 2440
rect 18414 2388 18420 2440
rect 18472 2388 18478 2440
rect 18800 2437 18828 2468
rect 19058 2456 19064 2508
rect 19116 2496 19122 2508
rect 19116 2468 19288 2496
rect 19116 2456 19122 2468
rect 19260 2437 19288 2468
rect 19426 2456 19432 2508
rect 19484 2496 19490 2508
rect 19484 2468 20392 2496
rect 19484 2456 19490 2468
rect 18785 2431 18843 2437
rect 18785 2397 18797 2431
rect 18831 2397 18843 2431
rect 18785 2391 18843 2397
rect 19245 2431 19303 2437
rect 19245 2397 19257 2431
rect 19291 2397 19303 2431
rect 19245 2391 19303 2397
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 19392 2400 19625 2428
rect 19392 2388 19398 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 19613 2391 19671 2397
rect 19978 2388 19984 2440
rect 20036 2388 20042 2440
rect 20364 2437 20392 2468
rect 21266 2456 21272 2508
rect 21324 2496 21330 2508
rect 22112 2496 22140 2604
rect 22646 2592 22652 2644
rect 22704 2632 22710 2644
rect 23753 2635 23811 2641
rect 23753 2632 23765 2635
rect 22704 2604 23765 2632
rect 22704 2592 22710 2604
rect 23753 2601 23765 2604
rect 23799 2601 23811 2635
rect 23753 2595 23811 2601
rect 24210 2592 24216 2644
rect 24268 2632 24274 2644
rect 25593 2635 25651 2641
rect 25593 2632 25605 2635
rect 24268 2604 25605 2632
rect 24268 2592 24274 2604
rect 25593 2601 25605 2604
rect 25639 2601 25651 2635
rect 25593 2595 25651 2601
rect 25866 2592 25872 2644
rect 25924 2632 25930 2644
rect 25924 2604 32720 2632
rect 25924 2592 25930 2604
rect 22186 2524 22192 2576
rect 22244 2564 22250 2576
rect 23385 2567 23443 2573
rect 23385 2564 23397 2567
rect 22244 2536 23397 2564
rect 22244 2524 22250 2536
rect 23385 2533 23397 2536
rect 23431 2533 23443 2567
rect 23385 2527 23443 2533
rect 23474 2524 23480 2576
rect 23532 2564 23538 2576
rect 24857 2567 24915 2573
rect 24857 2564 24869 2567
rect 23532 2536 24869 2564
rect 23532 2524 23538 2536
rect 24857 2533 24869 2536
rect 24903 2533 24915 2567
rect 25225 2567 25283 2573
rect 25225 2564 25237 2567
rect 24857 2527 24915 2533
rect 24964 2536 25237 2564
rect 21324 2468 21956 2496
rect 22112 2468 22876 2496
rect 21324 2456 21330 2468
rect 20349 2431 20407 2437
rect 20349 2397 20361 2431
rect 20395 2397 20407 2431
rect 20349 2391 20407 2397
rect 20717 2431 20775 2437
rect 20717 2397 20729 2431
rect 20763 2428 20775 2431
rect 20806 2428 20812 2440
rect 20763 2400 20812 2428
rect 20763 2397 20775 2400
rect 20717 2391 20775 2397
rect 20806 2388 20812 2400
rect 20864 2388 20870 2440
rect 21085 2431 21143 2437
rect 21085 2397 21097 2431
rect 21131 2397 21143 2431
rect 21085 2391 21143 2397
rect 15930 2360 15936 2372
rect 4212 2332 15148 2360
rect 15304 2332 15936 2360
rect 4212 2320 4218 2332
rect 10226 2252 10232 2304
rect 10284 2292 10290 2304
rect 13078 2292 13084 2304
rect 10284 2264 13084 2292
rect 10284 2252 10290 2264
rect 13078 2252 13084 2264
rect 13136 2252 13142 2304
rect 15304 2301 15332 2332
rect 15930 2320 15936 2332
rect 15988 2320 15994 2372
rect 19058 2320 19064 2372
rect 19116 2360 19122 2372
rect 19116 2332 20208 2360
rect 19116 2320 19122 2332
rect 15289 2295 15347 2301
rect 15289 2261 15301 2295
rect 15335 2261 15347 2295
rect 15289 2255 15347 2261
rect 15657 2295 15715 2301
rect 15657 2261 15669 2295
rect 15703 2292 15715 2295
rect 16298 2292 16304 2304
rect 15703 2264 16304 2292
rect 15703 2261 15715 2264
rect 15657 2255 15715 2261
rect 16298 2252 16304 2264
rect 16356 2252 16362 2304
rect 16393 2295 16451 2301
rect 16393 2261 16405 2295
rect 16439 2292 16451 2295
rect 16850 2292 16856 2304
rect 16439 2264 16856 2292
rect 16439 2261 16451 2264
rect 16393 2255 16451 2261
rect 16850 2252 16856 2264
rect 16908 2252 16914 2304
rect 17129 2295 17187 2301
rect 17129 2261 17141 2295
rect 17175 2292 17187 2295
rect 17218 2292 17224 2304
rect 17175 2264 17224 2292
rect 17175 2261 17187 2264
rect 17129 2255 17187 2261
rect 17218 2252 17224 2264
rect 17276 2252 17282 2304
rect 17497 2295 17555 2301
rect 17497 2261 17509 2295
rect 17543 2292 17555 2295
rect 17586 2292 17592 2304
rect 17543 2264 17592 2292
rect 17543 2261 17555 2264
rect 17497 2255 17555 2261
rect 17586 2252 17592 2264
rect 17644 2252 17650 2304
rect 17770 2252 17776 2304
rect 17828 2292 17834 2304
rect 17865 2295 17923 2301
rect 17865 2292 17877 2295
rect 17828 2264 17877 2292
rect 17828 2252 17834 2264
rect 17865 2261 17877 2264
rect 17911 2261 17923 2295
rect 17865 2255 17923 2261
rect 17954 2252 17960 2304
rect 18012 2292 18018 2304
rect 18233 2295 18291 2301
rect 18233 2292 18245 2295
rect 18012 2264 18245 2292
rect 18012 2252 18018 2264
rect 18233 2261 18245 2264
rect 18279 2261 18291 2295
rect 18233 2255 18291 2261
rect 18322 2252 18328 2304
rect 18380 2292 18386 2304
rect 18601 2295 18659 2301
rect 18601 2292 18613 2295
rect 18380 2264 18613 2292
rect 18380 2252 18386 2264
rect 18601 2261 18613 2264
rect 18647 2261 18659 2295
rect 18601 2255 18659 2261
rect 18690 2252 18696 2304
rect 18748 2292 18754 2304
rect 20180 2301 20208 2332
rect 20438 2320 20444 2372
rect 20496 2360 20502 2372
rect 21100 2360 21128 2391
rect 21726 2388 21732 2440
rect 21784 2428 21790 2440
rect 21821 2431 21879 2437
rect 21821 2428 21833 2431
rect 21784 2400 21833 2428
rect 21784 2388 21790 2400
rect 21821 2397 21833 2400
rect 21867 2397 21879 2431
rect 21928 2428 21956 2468
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 21928 2400 22201 2428
rect 21821 2391 21879 2397
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 22189 2391 22247 2397
rect 22554 2388 22560 2440
rect 22612 2388 22618 2440
rect 20496 2332 21128 2360
rect 20496 2320 20502 2332
rect 21450 2320 21456 2372
rect 21508 2360 21514 2372
rect 21508 2332 22784 2360
rect 21508 2320 21514 2332
rect 19797 2295 19855 2301
rect 19797 2292 19809 2295
rect 18748 2264 19809 2292
rect 18748 2252 18754 2264
rect 19797 2261 19809 2264
rect 19843 2261 19855 2295
rect 19797 2255 19855 2261
rect 20165 2295 20223 2301
rect 20165 2261 20177 2295
rect 20211 2261 20223 2295
rect 20165 2255 20223 2261
rect 20254 2252 20260 2304
rect 20312 2292 20318 2304
rect 20901 2295 20959 2301
rect 20901 2292 20913 2295
rect 20312 2264 20913 2292
rect 20312 2252 20318 2264
rect 20901 2261 20913 2264
rect 20947 2261 20959 2295
rect 20901 2255 20959 2261
rect 20990 2252 20996 2304
rect 21048 2292 21054 2304
rect 21542 2292 21548 2304
rect 21048 2264 21548 2292
rect 21048 2252 21054 2264
rect 21542 2252 21548 2264
rect 21600 2252 21606 2304
rect 21726 2252 21732 2304
rect 21784 2292 21790 2304
rect 22756 2301 22784 2332
rect 22373 2295 22431 2301
rect 22373 2292 22385 2295
rect 21784 2264 22385 2292
rect 21784 2252 21790 2264
rect 22373 2261 22385 2264
rect 22419 2261 22431 2295
rect 22373 2255 22431 2261
rect 22741 2295 22799 2301
rect 22741 2261 22753 2295
rect 22787 2261 22799 2295
rect 22848 2292 22876 2468
rect 22925 2431 22983 2437
rect 22925 2397 22937 2431
rect 22971 2428 22983 2431
rect 23014 2428 23020 2440
rect 22971 2400 23020 2428
rect 22971 2397 22983 2400
rect 22925 2391 22983 2397
rect 23014 2388 23020 2400
rect 23072 2388 23078 2440
rect 23566 2388 23572 2440
rect 23624 2388 23630 2440
rect 23934 2388 23940 2440
rect 23992 2388 23998 2440
rect 24486 2388 24492 2440
rect 24544 2428 24550 2440
rect 24673 2431 24731 2437
rect 24673 2428 24685 2431
rect 24544 2400 24685 2428
rect 24544 2388 24550 2400
rect 24673 2397 24685 2400
rect 24719 2397 24731 2431
rect 24673 2391 24731 2397
rect 23842 2320 23848 2372
rect 23900 2360 23906 2372
rect 24964 2360 24992 2536
rect 25225 2533 25237 2536
rect 25271 2533 25283 2567
rect 27798 2564 27804 2576
rect 25225 2527 25283 2533
rect 25424 2536 27804 2564
rect 25041 2431 25099 2437
rect 25041 2397 25053 2431
rect 25087 2428 25099 2431
rect 25314 2428 25320 2440
rect 25087 2400 25320 2428
rect 25087 2397 25099 2400
rect 25041 2391 25099 2397
rect 25314 2388 25320 2400
rect 25372 2388 25378 2440
rect 25424 2437 25452 2536
rect 27798 2524 27804 2536
rect 27856 2524 27862 2576
rect 26786 2496 26792 2508
rect 25792 2468 26792 2496
rect 25792 2437 25820 2468
rect 26786 2456 26792 2468
rect 26844 2456 26850 2508
rect 25409 2431 25467 2437
rect 25409 2397 25421 2431
rect 25455 2397 25467 2431
rect 25409 2391 25467 2397
rect 25777 2431 25835 2437
rect 25777 2397 25789 2431
rect 25823 2397 25835 2431
rect 25777 2391 25835 2397
rect 26145 2431 26203 2437
rect 26145 2397 26157 2431
rect 26191 2428 26203 2431
rect 26694 2428 26700 2440
rect 26191 2400 26700 2428
rect 26191 2397 26203 2400
rect 26145 2391 26203 2397
rect 26694 2388 26700 2400
rect 26752 2388 26758 2440
rect 30926 2388 30932 2440
rect 30984 2388 30990 2440
rect 31294 2388 31300 2440
rect 31352 2388 31358 2440
rect 31662 2388 31668 2440
rect 31720 2388 31726 2440
rect 32306 2388 32312 2440
rect 32364 2388 32370 2440
rect 32692 2437 32720 2604
rect 32858 2524 32864 2576
rect 32916 2524 32922 2576
rect 32677 2431 32735 2437
rect 32677 2397 32689 2431
rect 32723 2397 32735 2431
rect 32677 2391 32735 2397
rect 23900 2332 24992 2360
rect 23900 2320 23906 2332
rect 23109 2295 23167 2301
rect 23109 2292 23121 2295
rect 22848 2264 23121 2292
rect 22741 2255 22799 2261
rect 23109 2261 23121 2264
rect 23155 2261 23167 2295
rect 23109 2255 23167 2261
rect 23198 2252 23204 2304
rect 23256 2292 23262 2304
rect 24489 2295 24547 2301
rect 24489 2292 24501 2295
rect 23256 2264 24501 2292
rect 23256 2252 23262 2264
rect 24489 2261 24501 2264
rect 24535 2261 24547 2295
rect 24489 2255 24547 2261
rect 24578 2252 24584 2304
rect 24636 2292 24642 2304
rect 25961 2295 26019 2301
rect 25961 2292 25973 2295
rect 24636 2264 25973 2292
rect 24636 2252 24642 2264
rect 25961 2261 25973 2264
rect 26007 2261 26019 2295
rect 25961 2255 26019 2261
rect 31110 2252 31116 2304
rect 31168 2252 31174 2304
rect 31478 2252 31484 2304
rect 31536 2252 31542 2304
rect 31846 2252 31852 2304
rect 31904 2252 31910 2304
rect 32493 2295 32551 2301
rect 32493 2261 32505 2295
rect 32539 2292 32551 2295
rect 33410 2292 33416 2304
rect 32539 2264 33416 2292
rect 32539 2261 32551 2264
rect 32493 2255 32551 2261
rect 33410 2252 33416 2264
rect 33468 2252 33474 2304
rect 1104 2202 33324 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 9010 2202
rect 9062 2150 9074 2202
rect 9126 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 15010 2202
rect 15062 2150 15074 2202
rect 15126 2150 15138 2202
rect 15190 2150 15202 2202
rect 15254 2150 15266 2202
rect 15318 2150 21010 2202
rect 21062 2150 21074 2202
rect 21126 2150 21138 2202
rect 21190 2150 21202 2202
rect 21254 2150 21266 2202
rect 21318 2150 27010 2202
rect 27062 2150 27074 2202
rect 27126 2150 27138 2202
rect 27190 2150 27202 2202
rect 27254 2150 27266 2202
rect 27318 2150 33010 2202
rect 33062 2150 33074 2202
rect 33126 2150 33138 2202
rect 33190 2150 33202 2202
rect 33254 2150 33266 2202
rect 33318 2150 33324 2202
rect 1104 2128 33324 2150
rect 11054 2048 11060 2100
rect 11112 2088 11118 2100
rect 16206 2088 16212 2100
rect 11112 2060 16212 2088
rect 11112 2048 11118 2060
rect 16206 2048 16212 2060
rect 16264 2048 16270 2100
rect 16390 2048 16396 2100
rect 16448 2088 16454 2100
rect 19978 2088 19984 2100
rect 16448 2060 19984 2088
rect 16448 2048 16454 2060
rect 19978 2048 19984 2060
rect 20036 2048 20042 2100
rect 22370 2048 22376 2100
rect 22428 2088 22434 2100
rect 22428 2060 22692 2088
rect 22428 2048 22434 2060
rect 7466 1980 7472 2032
rect 7524 2020 7530 2032
rect 18414 2020 18420 2032
rect 7524 1992 18420 2020
rect 7524 1980 7530 1992
rect 18414 1980 18420 1992
rect 18472 1980 18478 2032
rect 18598 1980 18604 2032
rect 18656 2020 18662 2032
rect 22554 2020 22560 2032
rect 18656 1992 22560 2020
rect 18656 1980 18662 1992
rect 22554 1980 22560 1992
rect 22612 1980 22618 2032
rect 22664 2020 22692 2060
rect 23566 2048 23572 2100
rect 23624 2088 23630 2100
rect 28166 2088 28172 2100
rect 23624 2060 28172 2088
rect 23624 2048 23630 2060
rect 28166 2048 28172 2060
rect 28224 2048 28230 2100
rect 31294 2020 31300 2032
rect 22664 1992 31300 2020
rect 31294 1980 31300 1992
rect 31352 1980 31358 2032
rect 17126 1912 17132 1964
rect 17184 1952 17190 1964
rect 20438 1952 20444 1964
rect 17184 1924 20444 1952
rect 17184 1912 17190 1924
rect 20438 1912 20444 1924
rect 20496 1912 20502 1964
rect 22094 1912 22100 1964
rect 22152 1952 22158 1964
rect 30926 1952 30932 1964
rect 22152 1924 30932 1952
rect 22152 1912 22158 1924
rect 30926 1912 30932 1924
rect 30984 1912 30990 1964
rect 7190 1844 7196 1896
rect 7248 1884 7254 1896
rect 17310 1884 17316 1896
rect 7248 1856 17316 1884
rect 7248 1844 7254 1856
rect 17310 1844 17316 1856
rect 17368 1844 17374 1896
rect 19150 1844 19156 1896
rect 19208 1884 19214 1896
rect 31662 1884 31668 1896
rect 19208 1856 31668 1884
rect 19208 1844 19214 1856
rect 31662 1844 31668 1856
rect 31720 1844 31726 1896
rect 8294 1776 8300 1828
rect 8352 1816 8358 1828
rect 19334 1816 19340 1828
rect 8352 1788 19340 1816
rect 8352 1776 8358 1788
rect 19334 1776 19340 1788
rect 19392 1776 19398 1828
rect 24302 1776 24308 1828
rect 24360 1816 24366 1828
rect 27706 1816 27712 1828
rect 24360 1788 27712 1816
rect 24360 1776 24366 1788
rect 27706 1776 27712 1788
rect 27764 1776 27770 1828
rect 7374 1708 7380 1760
rect 7432 1748 7438 1760
rect 18046 1748 18052 1760
rect 7432 1720 18052 1748
rect 7432 1708 7438 1720
rect 18046 1708 18052 1720
rect 18104 1708 18110 1760
rect 4430 1640 4436 1692
rect 4488 1680 4494 1692
rect 16942 1680 16948 1692
rect 4488 1652 16948 1680
rect 4488 1640 4494 1652
rect 16942 1640 16948 1652
rect 17000 1640 17006 1692
rect 29178 1680 29184 1692
rect 22066 1652 29184 1680
rect 14458 1572 14464 1624
rect 14516 1612 14522 1624
rect 22066 1612 22094 1652
rect 29178 1640 29184 1652
rect 29236 1640 29242 1692
rect 14516 1584 22094 1612
rect 14516 1572 14522 1584
rect 27338 1572 27344 1624
rect 27396 1612 27402 1624
rect 29638 1612 29644 1624
rect 27396 1584 29644 1612
rect 27396 1572 27402 1584
rect 29638 1572 29644 1584
rect 29696 1572 29702 1624
rect 15654 1504 15660 1556
rect 15712 1544 15718 1556
rect 23014 1544 23020 1556
rect 15712 1516 23020 1544
rect 15712 1504 15718 1516
rect 23014 1504 23020 1516
rect 23072 1504 23078 1556
rect 28442 1504 28448 1556
rect 28500 1544 28506 1556
rect 30834 1544 30840 1556
rect 28500 1516 30840 1544
rect 28500 1504 28506 1516
rect 30834 1504 30840 1516
rect 30892 1504 30898 1556
rect 14642 1436 14648 1488
rect 14700 1476 14706 1488
rect 18598 1476 18604 1488
rect 14700 1448 18604 1476
rect 14700 1436 14706 1448
rect 18598 1436 18604 1448
rect 18656 1436 18662 1488
rect 19518 1436 19524 1488
rect 19576 1476 19582 1488
rect 19886 1476 19892 1488
rect 19576 1448 19892 1476
rect 19576 1436 19582 1448
rect 19886 1436 19892 1448
rect 19944 1436 19950 1488
rect 21542 1436 21548 1488
rect 21600 1476 21606 1488
rect 32306 1476 32312 1488
rect 21600 1448 32312 1476
rect 21600 1436 21606 1448
rect 32306 1436 32312 1448
rect 32364 1436 32370 1488
rect 19702 1368 19708 1420
rect 19760 1408 19766 1420
rect 20254 1408 20260 1420
rect 19760 1380 20260 1408
rect 19760 1368 19766 1380
rect 20254 1368 20260 1380
rect 20312 1368 20318 1420
rect 21082 1368 21088 1420
rect 21140 1408 21146 1420
rect 21726 1408 21732 1420
rect 21140 1380 21732 1408
rect 21140 1368 21146 1380
rect 21726 1368 21732 1380
rect 21784 1368 21790 1420
rect 27154 1368 27160 1420
rect 27212 1408 27218 1420
rect 27614 1408 27620 1420
rect 27212 1380 27620 1408
rect 27212 1368 27218 1380
rect 27614 1368 27620 1380
rect 27672 1368 27678 1420
rect 28258 1368 28264 1420
rect 28316 1408 28322 1420
rect 29914 1408 29920 1420
rect 28316 1380 29920 1408
rect 28316 1368 28322 1380
rect 29914 1368 29920 1380
rect 29972 1368 29978 1420
rect 9306 1300 9312 1352
rect 9364 1340 9370 1352
rect 14550 1340 14556 1352
rect 9364 1312 14556 1340
rect 9364 1300 9370 1312
rect 14550 1300 14556 1312
rect 14608 1300 14614 1352
rect 9490 1232 9496 1284
rect 9548 1272 9554 1284
rect 15838 1272 15844 1284
rect 9548 1244 15844 1272
rect 9548 1232 9554 1244
rect 15838 1232 15844 1244
rect 15896 1232 15902 1284
rect 14918 688 14924 740
rect 14976 728 14982 740
rect 25498 728 25504 740
rect 14976 700 25504 728
rect 14976 688 14982 700
rect 25498 688 25504 700
rect 25556 688 25562 740
rect 14826 484 14832 536
rect 14884 524 14890 536
rect 28534 524 28540 536
rect 14884 496 28540 524
rect 14884 484 14890 496
rect 28534 484 28540 496
rect 28592 484 28598 536
rect 14366 416 14372 468
rect 14424 456 14430 468
rect 28350 456 28356 468
rect 14424 428 28356 456
rect 14424 416 14430 428
rect 28350 416 28356 428
rect 28408 416 28414 468
rect 12250 348 12256 400
rect 12308 388 12314 400
rect 26510 388 26516 400
rect 12308 360 26516 388
rect 12308 348 12314 360
rect 26510 348 26516 360
rect 26568 348 26574 400
rect 13170 280 13176 332
rect 13228 320 13234 332
rect 28718 320 28724 332
rect 13228 292 28724 320
rect 13228 280 13234 292
rect 28718 280 28724 292
rect 28776 280 28782 332
rect 12618 212 12624 264
rect 12676 252 12682 264
rect 12676 224 13308 252
rect 12676 212 12682 224
rect 12802 144 12808 196
rect 12860 184 12866 196
rect 13280 184 13308 224
rect 15010 212 15016 264
rect 15068 252 15074 264
rect 29546 252 29552 264
rect 15068 224 29552 252
rect 15068 212 15074 224
rect 29546 212 29552 224
rect 29604 212 29610 264
rect 27246 184 27252 196
rect 12860 156 13216 184
rect 13280 156 27252 184
rect 12860 144 12866 156
rect 13078 76 13084 128
rect 13136 76 13142 128
rect 13188 116 13216 156
rect 27246 144 27252 156
rect 27304 144 27310 196
rect 27430 116 27436 128
rect 13188 88 27436 116
rect 27430 76 27436 88
rect 27488 76 27494 128
rect 27798 76 27804 128
rect 27856 76 27862 128
rect 13096 48 13124 76
rect 27816 48 27844 76
rect 13096 20 27844 48
<< via1 >>
rect 14372 9052 14424 9104
rect 25780 9052 25832 9104
rect 12808 8984 12860 9036
rect 28540 8984 28592 9036
rect 17316 8916 17368 8968
rect 30932 8916 30984 8968
rect 11244 8848 11296 8900
rect 28264 8848 28316 8900
rect 8024 8780 8076 8832
rect 14832 8780 14884 8832
rect 20628 8780 20680 8832
rect 27436 8780 27488 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 9010 8678 9062 8730
rect 9074 8678 9126 8730
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 15010 8678 15062 8730
rect 15074 8678 15126 8730
rect 15138 8678 15190 8730
rect 15202 8678 15254 8730
rect 15266 8678 15318 8730
rect 21010 8678 21062 8730
rect 21074 8678 21126 8730
rect 21138 8678 21190 8730
rect 21202 8678 21254 8730
rect 21266 8678 21318 8730
rect 27010 8678 27062 8730
rect 27074 8678 27126 8730
rect 27138 8678 27190 8730
rect 27202 8678 27254 8730
rect 27266 8678 27318 8730
rect 33010 8678 33062 8730
rect 33074 8678 33126 8730
rect 33138 8678 33190 8730
rect 33202 8678 33254 8730
rect 33266 8678 33318 8730
rect 1492 8576 1544 8628
rect 2872 8576 2924 8628
rect 4620 8576 4672 8628
rect 6184 8576 6236 8628
rect 7748 8576 7800 8628
rect 9404 8576 9456 8628
rect 12440 8576 12492 8628
rect 14004 8576 14056 8628
rect 15568 8576 15620 8628
rect 17132 8576 17184 8628
rect 18696 8576 18748 8628
rect 11060 8508 11112 8560
rect 19708 8576 19760 8628
rect 20260 8576 20312 8628
rect 21824 8576 21876 8628
rect 23388 8576 23440 8628
rect 24952 8576 25004 8628
rect 26516 8576 26568 8628
rect 28080 8576 28132 8628
rect 29644 8576 29696 8628
rect 31116 8619 31168 8628
rect 31116 8585 31125 8619
rect 31125 8585 31159 8619
rect 31159 8585 31168 8619
rect 31116 8576 31168 8585
rect 31208 8576 31260 8628
rect 32772 8576 32824 8628
rect 8024 8440 8076 8492
rect 11244 8483 11296 8492
rect 11244 8449 11253 8483
rect 11253 8449 11287 8483
rect 11287 8449 11296 8483
rect 11244 8440 11296 8449
rect 12808 8483 12860 8492
rect 12808 8449 12817 8483
rect 12817 8449 12851 8483
rect 12851 8449 12860 8483
rect 12808 8440 12860 8449
rect 14372 8483 14424 8492
rect 14372 8449 14381 8483
rect 14381 8449 14415 8483
rect 14415 8449 14424 8483
rect 14372 8440 14424 8449
rect 17408 8440 17460 8492
rect 25320 8508 25372 8560
rect 30656 8508 30708 8560
rect 20628 8483 20680 8492
rect 20628 8449 20637 8483
rect 20637 8449 20671 8483
rect 20671 8449 20680 8483
rect 20628 8440 20680 8449
rect 24860 8440 24912 8492
rect 27988 8440 28040 8492
rect 28724 8440 28776 8492
rect 29736 8483 29788 8492
rect 29736 8449 29745 8483
rect 29745 8449 29779 8483
rect 29779 8449 29788 8483
rect 29736 8440 29788 8449
rect 30932 8483 30984 8492
rect 30932 8449 30941 8483
rect 30941 8449 30975 8483
rect 30975 8449 30984 8483
rect 30932 8440 30984 8449
rect 31300 8483 31352 8492
rect 31300 8449 31309 8483
rect 31309 8449 31343 8483
rect 31343 8449 31352 8483
rect 31300 8440 31352 8449
rect 5540 8236 5592 8288
rect 9496 8236 9548 8288
rect 10876 8304 10928 8356
rect 13820 8304 13872 8356
rect 17408 8304 17460 8356
rect 19432 8304 19484 8356
rect 30840 8372 30892 8424
rect 31024 8372 31076 8424
rect 32404 8440 32456 8492
rect 29460 8304 29512 8356
rect 33048 8304 33100 8356
rect 24768 8236 24820 8288
rect 32496 8279 32548 8288
rect 32496 8245 32505 8279
rect 32505 8245 32539 8279
rect 32539 8245 32548 8279
rect 32496 8236 32548 8245
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 13950 8134 14002 8186
rect 14014 8134 14066 8186
rect 14078 8134 14130 8186
rect 14142 8134 14194 8186
rect 14206 8134 14258 8186
rect 19950 8134 20002 8186
rect 20014 8134 20066 8186
rect 20078 8134 20130 8186
rect 20142 8134 20194 8186
rect 20206 8134 20258 8186
rect 25950 8134 26002 8186
rect 26014 8134 26066 8186
rect 26078 8134 26130 8186
rect 26142 8134 26194 8186
rect 26206 8134 26258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 17224 8032 17276 8084
rect 24952 8032 25004 8084
rect 31392 8075 31444 8084
rect 31392 8041 31401 8075
rect 31401 8041 31435 8075
rect 31435 8041 31444 8075
rect 31392 8032 31444 8041
rect 31760 8075 31812 8084
rect 31760 8041 31769 8075
rect 31769 8041 31803 8075
rect 31803 8041 31812 8075
rect 31760 8032 31812 8041
rect 32312 8032 32364 8084
rect 16580 7964 16632 8016
rect 1124 7896 1176 7948
rect 24216 7896 24268 7948
rect 24584 7896 24636 7948
rect 14372 7828 14424 7880
rect 23020 7828 23072 7880
rect 31208 7871 31260 7880
rect 31208 7837 31217 7871
rect 31217 7837 31251 7871
rect 31251 7837 31260 7871
rect 31208 7828 31260 7837
rect 31668 7828 31720 7880
rect 1400 7692 1452 7744
rect 17592 7760 17644 7812
rect 19156 7760 19208 7812
rect 12348 7692 12400 7744
rect 19340 7692 19392 7744
rect 32496 7735 32548 7744
rect 32496 7701 32505 7735
rect 32505 7701 32539 7735
rect 32539 7701 32548 7735
rect 32496 7692 32548 7701
rect 33600 7692 33652 7744
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 9010 7590 9062 7642
rect 9074 7590 9126 7642
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 15010 7590 15062 7642
rect 15074 7590 15126 7642
rect 15138 7590 15190 7642
rect 15202 7590 15254 7642
rect 15266 7590 15318 7642
rect 21010 7590 21062 7642
rect 21074 7590 21126 7642
rect 21138 7590 21190 7642
rect 21202 7590 21254 7642
rect 21266 7590 21318 7642
rect 27010 7590 27062 7642
rect 27074 7590 27126 7642
rect 27138 7590 27190 7642
rect 27202 7590 27254 7642
rect 27266 7590 27318 7642
rect 33010 7590 33062 7642
rect 33074 7590 33126 7642
rect 33138 7590 33190 7642
rect 33202 7590 33254 7642
rect 33266 7590 33318 7642
rect 5540 7488 5592 7540
rect 11060 7531 11112 7540
rect 11060 7497 11069 7531
rect 11069 7497 11103 7531
rect 11103 7497 11112 7531
rect 11060 7488 11112 7497
rect 13820 7488 13872 7540
rect 14832 7531 14884 7540
rect 14832 7497 14841 7531
rect 14841 7497 14875 7531
rect 14875 7497 14884 7531
rect 14832 7488 14884 7497
rect 17592 7531 17644 7540
rect 17592 7497 17601 7531
rect 17601 7497 17635 7531
rect 17635 7497 17644 7531
rect 17592 7488 17644 7497
rect 24124 7488 24176 7540
rect 24768 7531 24820 7540
rect 24768 7497 24777 7531
rect 24777 7497 24811 7531
rect 24811 7497 24820 7531
rect 24768 7488 24820 7497
rect 25320 7531 25372 7540
rect 25320 7497 25329 7531
rect 25329 7497 25363 7531
rect 25363 7497 25372 7531
rect 25320 7488 25372 7497
rect 27436 7488 27488 7540
rect 27988 7531 28040 7540
rect 27988 7497 27997 7531
rect 27997 7497 28031 7531
rect 28031 7497 28040 7531
rect 27988 7488 28040 7497
rect 28264 7531 28316 7540
rect 28264 7497 28273 7531
rect 28273 7497 28307 7531
rect 28307 7497 28316 7531
rect 28264 7488 28316 7497
rect 28540 7531 28592 7540
rect 28540 7497 28549 7531
rect 28549 7497 28583 7531
rect 28583 7497 28592 7531
rect 28540 7488 28592 7497
rect 29460 7531 29512 7540
rect 29460 7497 29469 7531
rect 29469 7497 29503 7531
rect 29503 7497 29512 7531
rect 29460 7488 29512 7497
rect 30840 7488 30892 7540
rect 33416 7488 33468 7540
rect 1216 7284 1268 7336
rect 9588 7352 9640 7404
rect 12348 7395 12400 7404
rect 12348 7361 12357 7395
rect 12357 7361 12391 7395
rect 12391 7361 12400 7395
rect 12348 7352 12400 7361
rect 14372 7395 14424 7404
rect 14372 7361 14381 7395
rect 14381 7361 14415 7395
rect 14415 7361 14424 7395
rect 14372 7352 14424 7361
rect 14924 7352 14976 7404
rect 18052 7395 18104 7404
rect 18052 7361 18061 7395
rect 18061 7361 18095 7395
rect 18095 7361 18104 7395
rect 18052 7352 18104 7361
rect 19800 7395 19852 7404
rect 19800 7361 19809 7395
rect 19809 7361 19843 7395
rect 19843 7361 19852 7395
rect 19800 7352 19852 7361
rect 21824 7395 21876 7404
rect 21824 7361 21833 7395
rect 21833 7361 21867 7395
rect 21867 7361 21876 7395
rect 21824 7352 21876 7361
rect 17224 7284 17276 7336
rect 26884 7420 26936 7472
rect 24216 7395 24268 7404
rect 24216 7361 24225 7395
rect 24225 7361 24259 7395
rect 24259 7361 24268 7395
rect 24216 7352 24268 7361
rect 1676 7216 1728 7268
rect 24768 7284 24820 7336
rect 9496 7148 9548 7200
rect 17960 7191 18012 7200
rect 17960 7157 17969 7191
rect 17969 7157 18003 7191
rect 18003 7157 18012 7191
rect 17960 7148 18012 7157
rect 18236 7191 18288 7200
rect 18236 7157 18245 7191
rect 18245 7157 18279 7191
rect 18279 7157 18288 7191
rect 18236 7148 18288 7157
rect 22008 7191 22060 7200
rect 22008 7157 22017 7191
rect 22017 7157 22051 7191
rect 22051 7157 22060 7191
rect 22008 7148 22060 7157
rect 22284 7191 22336 7200
rect 22284 7157 22293 7191
rect 22293 7157 22327 7191
rect 22327 7157 22336 7191
rect 22284 7148 22336 7157
rect 25596 7352 25648 7404
rect 27620 7352 27672 7404
rect 27988 7352 28040 7404
rect 28448 7395 28500 7404
rect 28448 7361 28457 7395
rect 28457 7361 28491 7395
rect 28491 7361 28500 7395
rect 28448 7352 28500 7361
rect 25688 7284 25740 7336
rect 26792 7284 26844 7336
rect 29644 7395 29696 7404
rect 29644 7361 29653 7395
rect 29653 7361 29687 7395
rect 29687 7361 29696 7395
rect 29644 7352 29696 7361
rect 30472 7352 30524 7404
rect 31392 7352 31444 7404
rect 30380 7284 30432 7336
rect 25872 7216 25924 7268
rect 30564 7148 30616 7200
rect 32864 7191 32916 7200
rect 32864 7157 32873 7191
rect 32873 7157 32907 7191
rect 32907 7157 32916 7191
rect 32864 7148 32916 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 13950 7046 14002 7098
rect 14014 7046 14066 7098
rect 14078 7046 14130 7098
rect 14142 7046 14194 7098
rect 14206 7046 14258 7098
rect 19950 7046 20002 7098
rect 20014 7046 20066 7098
rect 20078 7046 20130 7098
rect 20142 7046 20194 7098
rect 20206 7046 20258 7098
rect 25950 7046 26002 7098
rect 26014 7046 26066 7098
rect 26078 7046 26130 7098
rect 26142 7046 26194 7098
rect 26206 7046 26258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 848 6944 900 6996
rect 21824 6944 21876 6996
rect 24768 6944 24820 6996
rect 31852 6944 31904 6996
rect 2688 6876 2740 6928
rect 18052 6876 18104 6928
rect 1768 6808 1820 6860
rect 1308 6740 1360 6792
rect 16488 6808 16540 6860
rect 24124 6876 24176 6928
rect 30932 6876 30984 6928
rect 30380 6808 30432 6860
rect 16120 6604 16172 6656
rect 19800 6604 19852 6656
rect 20444 6647 20496 6656
rect 20444 6613 20453 6647
rect 20453 6613 20487 6647
rect 20487 6613 20496 6647
rect 20444 6604 20496 6613
rect 24492 6672 24544 6724
rect 24676 6783 24728 6792
rect 24676 6749 24685 6783
rect 24685 6749 24719 6783
rect 24719 6749 24728 6783
rect 24676 6740 24728 6749
rect 25412 6740 25464 6792
rect 26424 6740 26476 6792
rect 28080 6740 28132 6792
rect 31760 6740 31812 6792
rect 26608 6672 26660 6724
rect 26700 6672 26752 6724
rect 24400 6647 24452 6656
rect 24400 6613 24409 6647
rect 24409 6613 24443 6647
rect 24443 6613 24452 6647
rect 24400 6604 24452 6613
rect 24860 6647 24912 6656
rect 24860 6613 24869 6647
rect 24869 6613 24903 6647
rect 24903 6613 24912 6647
rect 24860 6604 24912 6613
rect 25136 6647 25188 6656
rect 25136 6613 25145 6647
rect 25145 6613 25179 6647
rect 25179 6613 25188 6647
rect 25136 6604 25188 6613
rect 25780 6604 25832 6656
rect 28724 6647 28776 6656
rect 28724 6613 28733 6647
rect 28733 6613 28767 6647
rect 28767 6613 28776 6647
rect 28724 6604 28776 6613
rect 33416 6672 33468 6724
rect 32864 6647 32916 6656
rect 32864 6613 32873 6647
rect 32873 6613 32907 6647
rect 32907 6613 32916 6647
rect 32864 6604 32916 6613
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 9010 6502 9062 6554
rect 9074 6502 9126 6554
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 15010 6502 15062 6554
rect 15074 6502 15126 6554
rect 15138 6502 15190 6554
rect 15202 6502 15254 6554
rect 15266 6502 15318 6554
rect 21010 6502 21062 6554
rect 21074 6502 21126 6554
rect 21138 6502 21190 6554
rect 21202 6502 21254 6554
rect 21266 6502 21318 6554
rect 27010 6502 27062 6554
rect 27074 6502 27126 6554
rect 27138 6502 27190 6554
rect 27202 6502 27254 6554
rect 27266 6502 27318 6554
rect 33010 6502 33062 6554
rect 33074 6502 33126 6554
rect 33138 6502 33190 6554
rect 33202 6502 33254 6554
rect 33266 6502 33318 6554
rect 2596 6400 2648 6452
rect 15568 6400 15620 6452
rect 15108 6332 15160 6384
rect 19156 6443 19208 6452
rect 19156 6409 19165 6443
rect 19165 6409 19199 6443
rect 19199 6409 19208 6443
rect 19156 6400 19208 6409
rect 19708 6400 19760 6452
rect 24400 6400 24452 6452
rect 24492 6400 24544 6452
rect 2780 6196 2832 6248
rect 16120 6196 16172 6248
rect 18972 6307 19024 6316
rect 18972 6273 18981 6307
rect 18981 6273 19015 6307
rect 19015 6273 19024 6307
rect 18972 6264 19024 6273
rect 19432 6332 19484 6384
rect 25136 6332 25188 6384
rect 29736 6443 29788 6452
rect 29736 6409 29745 6443
rect 29745 6409 29779 6443
rect 29779 6409 29788 6443
rect 29736 6400 29788 6409
rect 32864 6443 32916 6452
rect 32864 6409 32873 6443
rect 32873 6409 32907 6443
rect 32907 6409 32916 6443
rect 32864 6400 32916 6409
rect 31208 6332 31260 6384
rect 24584 6264 24636 6316
rect 29920 6307 29972 6316
rect 29920 6273 29929 6307
rect 29929 6273 29963 6307
rect 29963 6273 29972 6307
rect 29920 6264 29972 6273
rect 32312 6307 32364 6316
rect 32312 6273 32321 6307
rect 32321 6273 32355 6307
rect 32355 6273 32364 6307
rect 32312 6264 32364 6273
rect 31024 6196 31076 6248
rect 18972 6060 19024 6112
rect 32496 6103 32548 6112
rect 32496 6069 32505 6103
rect 32505 6069 32539 6103
rect 32539 6069 32548 6103
rect 32496 6060 32548 6069
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 13950 5958 14002 6010
rect 14014 5958 14066 6010
rect 14078 5958 14130 6010
rect 14142 5958 14194 6010
rect 14206 5958 14258 6010
rect 19950 5958 20002 6010
rect 20014 5958 20066 6010
rect 20078 5958 20130 6010
rect 20142 5958 20194 6010
rect 20206 5958 20258 6010
rect 25950 5958 26002 6010
rect 26014 5958 26066 6010
rect 26078 5958 26130 6010
rect 26142 5958 26194 6010
rect 26206 5958 26258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 17040 5899 17092 5908
rect 17040 5865 17049 5899
rect 17049 5865 17083 5899
rect 17083 5865 17092 5899
rect 17040 5856 17092 5865
rect 20444 5856 20496 5908
rect 30656 5856 30708 5908
rect 31300 5856 31352 5908
rect 9588 5788 9640 5840
rect 24860 5788 24912 5840
rect 32864 5831 32916 5840
rect 32864 5797 32873 5831
rect 32873 5797 32907 5831
rect 32907 5797 32916 5831
rect 32864 5788 32916 5797
rect 25872 5720 25924 5772
rect 17500 5695 17552 5704
rect 17500 5661 17509 5695
rect 17509 5661 17543 5695
rect 17543 5661 17552 5695
rect 17500 5652 17552 5661
rect 30840 5695 30892 5704
rect 30840 5661 30849 5695
rect 30849 5661 30883 5695
rect 30883 5661 30892 5695
rect 30840 5652 30892 5661
rect 30932 5652 30984 5704
rect 31668 5584 31720 5636
rect 31392 5516 31444 5568
rect 33416 5516 33468 5568
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 9010 5414 9062 5466
rect 9074 5414 9126 5466
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 15010 5414 15062 5466
rect 15074 5414 15126 5466
rect 15138 5414 15190 5466
rect 15202 5414 15254 5466
rect 15266 5414 15318 5466
rect 21010 5414 21062 5466
rect 21074 5414 21126 5466
rect 21138 5414 21190 5466
rect 21202 5414 21254 5466
rect 21266 5414 21318 5466
rect 27010 5414 27062 5466
rect 27074 5414 27126 5466
rect 27138 5414 27190 5466
rect 27202 5414 27254 5466
rect 27266 5414 27318 5466
rect 33010 5414 33062 5466
rect 33074 5414 33126 5466
rect 33138 5414 33190 5466
rect 33202 5414 33254 5466
rect 33266 5414 33318 5466
rect 3424 5244 3476 5296
rect 13452 5312 13504 5364
rect 15568 5355 15620 5364
rect 15568 5321 15577 5355
rect 15577 5321 15611 5355
rect 15611 5321 15620 5355
rect 15568 5312 15620 5321
rect 16396 5355 16448 5364
rect 16396 5321 16405 5355
rect 16405 5321 16439 5355
rect 16439 5321 16448 5355
rect 16396 5312 16448 5321
rect 32312 5312 32364 5364
rect 32864 5355 32916 5364
rect 32864 5321 32873 5355
rect 32873 5321 32907 5355
rect 32907 5321 32916 5355
rect 32864 5312 32916 5321
rect 7380 5244 7432 5296
rect 15200 5244 15252 5296
rect 15660 5244 15712 5296
rect 19432 5244 19484 5296
rect 3148 5176 3200 5228
rect 10048 5176 10100 5228
rect 13636 5176 13688 5228
rect 14740 5176 14792 5228
rect 16948 5176 17000 5228
rect 18236 5176 18288 5228
rect 28632 5176 28684 5228
rect 13268 5108 13320 5160
rect 15476 5040 15528 5092
rect 17316 5040 17368 5092
rect 17960 5108 18012 5160
rect 21732 5040 21784 5092
rect 32404 5040 32456 5092
rect 12072 4972 12124 5024
rect 17132 4972 17184 5024
rect 32496 5015 32548 5024
rect 32496 4981 32505 5015
rect 32505 4981 32539 5015
rect 32539 4981 32548 5015
rect 32496 4972 32548 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 13950 4870 14002 4922
rect 14014 4870 14066 4922
rect 14078 4870 14130 4922
rect 14142 4870 14194 4922
rect 14206 4870 14258 4922
rect 19950 4870 20002 4922
rect 20014 4870 20066 4922
rect 20078 4870 20130 4922
rect 20142 4870 20194 4922
rect 20206 4870 20258 4922
rect 25950 4870 26002 4922
rect 26014 4870 26066 4922
rect 26078 4870 26130 4922
rect 26142 4870 26194 4922
rect 26206 4870 26258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 3148 4811 3200 4820
rect 3148 4777 3157 4811
rect 3157 4777 3191 4811
rect 3191 4777 3200 4811
rect 3148 4768 3200 4777
rect 3424 4811 3476 4820
rect 3424 4777 3433 4811
rect 3433 4777 3467 4811
rect 3467 4777 3476 4811
rect 3424 4768 3476 4777
rect 7380 4811 7432 4820
rect 7380 4777 7389 4811
rect 7389 4777 7423 4811
rect 7423 4777 7432 4811
rect 7380 4768 7432 4777
rect 10968 4768 11020 4820
rect 6184 4632 6236 4684
rect 5816 4564 5868 4616
rect 8852 4564 8904 4616
rect 11704 4700 11756 4752
rect 11520 4632 11572 4684
rect 11336 4607 11388 4616
rect 11336 4573 11345 4607
rect 11345 4573 11379 4607
rect 11379 4573 11388 4607
rect 11336 4564 11388 4573
rect 12072 4811 12124 4820
rect 12072 4777 12081 4811
rect 12081 4777 12115 4811
rect 12115 4777 12124 4811
rect 12072 4768 12124 4777
rect 13268 4743 13320 4752
rect 13268 4709 13277 4743
rect 13277 4709 13311 4743
rect 13311 4709 13320 4743
rect 13268 4700 13320 4709
rect 11980 4632 12032 4684
rect 15384 4811 15436 4820
rect 15384 4777 15393 4811
rect 15393 4777 15427 4811
rect 15427 4777 15436 4811
rect 15384 4768 15436 4777
rect 15936 4811 15988 4820
rect 15936 4777 15945 4811
rect 15945 4777 15979 4811
rect 15979 4777 15988 4811
rect 15936 4768 15988 4777
rect 16212 4811 16264 4820
rect 16212 4777 16221 4811
rect 16221 4777 16255 4811
rect 16255 4777 16264 4811
rect 16212 4768 16264 4777
rect 22008 4768 22060 4820
rect 16396 4700 16448 4752
rect 6000 4496 6052 4548
rect 11152 4496 11204 4548
rect 12256 4607 12308 4616
rect 12256 4573 12265 4607
rect 12265 4573 12299 4607
rect 12299 4573 12308 4607
rect 12256 4564 12308 4573
rect 12532 4607 12584 4616
rect 12532 4573 12541 4607
rect 12541 4573 12575 4607
rect 12575 4573 12584 4607
rect 12532 4564 12584 4573
rect 13084 4607 13136 4616
rect 13084 4573 13093 4607
rect 13093 4573 13127 4607
rect 13127 4573 13136 4607
rect 13084 4564 13136 4573
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 13636 4607 13688 4616
rect 13636 4573 13645 4607
rect 13645 4573 13679 4607
rect 13679 4573 13688 4607
rect 13636 4564 13688 4573
rect 20628 4632 20680 4684
rect 23204 4700 23256 4752
rect 31760 4632 31812 4684
rect 12072 4496 12124 4548
rect 15752 4607 15804 4616
rect 15752 4573 15761 4607
rect 15761 4573 15795 4607
rect 15795 4573 15804 4607
rect 15752 4564 15804 4573
rect 25136 4564 25188 4616
rect 27804 4564 27856 4616
rect 27896 4607 27948 4616
rect 27896 4573 27905 4607
rect 27905 4573 27939 4607
rect 27939 4573 27948 4607
rect 27896 4564 27948 4573
rect 28264 4607 28316 4616
rect 28264 4573 28273 4607
rect 28273 4573 28307 4607
rect 28307 4573 28316 4607
rect 28264 4564 28316 4573
rect 10140 4428 10192 4480
rect 11060 4428 11112 4480
rect 11244 4471 11296 4480
rect 11244 4437 11253 4471
rect 11253 4437 11287 4471
rect 11287 4437 11296 4471
rect 11244 4428 11296 4437
rect 11612 4428 11664 4480
rect 11796 4471 11848 4480
rect 11796 4437 11805 4471
rect 11805 4437 11839 4471
rect 11839 4437 11848 4471
rect 11796 4428 11848 4437
rect 12440 4471 12492 4480
rect 12440 4437 12449 4471
rect 12449 4437 12483 4471
rect 12483 4437 12492 4471
rect 12440 4428 12492 4437
rect 12716 4471 12768 4480
rect 12716 4437 12725 4471
rect 12725 4437 12759 4471
rect 12759 4437 12768 4471
rect 12716 4428 12768 4437
rect 14832 4428 14884 4480
rect 19248 4496 19300 4548
rect 27528 4496 27580 4548
rect 31852 4564 31904 4616
rect 32864 4743 32916 4752
rect 32864 4709 32873 4743
rect 32873 4709 32907 4743
rect 32907 4709 32916 4743
rect 32864 4700 32916 4709
rect 15200 4428 15252 4480
rect 15568 4428 15620 4480
rect 16488 4428 16540 4480
rect 24492 4428 24544 4480
rect 27804 4428 27856 4480
rect 33416 4428 33468 4480
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 9010 4326 9062 4378
rect 9074 4326 9126 4378
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 15010 4326 15062 4378
rect 15074 4326 15126 4378
rect 15138 4326 15190 4378
rect 15202 4326 15254 4378
rect 15266 4326 15318 4378
rect 21010 4326 21062 4378
rect 21074 4326 21126 4378
rect 21138 4326 21190 4378
rect 21202 4326 21254 4378
rect 21266 4326 21318 4378
rect 27010 4326 27062 4378
rect 27074 4326 27126 4378
rect 27138 4326 27190 4378
rect 27202 4326 27254 4378
rect 27266 4326 27318 4378
rect 33010 4326 33062 4378
rect 33074 4326 33126 4378
rect 33138 4326 33190 4378
rect 33202 4326 33254 4378
rect 33266 4326 33318 4378
rect 2688 4267 2740 4276
rect 2688 4233 2697 4267
rect 2697 4233 2731 4267
rect 2731 4233 2740 4267
rect 2688 4224 2740 4233
rect 2412 4088 2464 4140
rect 2596 4088 2648 4140
rect 2872 4020 2924 4072
rect 2780 3952 2832 4004
rect 7012 4267 7064 4276
rect 7012 4233 7021 4267
rect 7021 4233 7055 4267
rect 7055 4233 7064 4267
rect 7012 4224 7064 4233
rect 10784 4224 10836 4276
rect 12256 4224 12308 4276
rect 12440 4224 12492 4276
rect 20444 4224 20496 4276
rect 3424 4131 3476 4140
rect 3424 4097 3433 4131
rect 3433 4097 3467 4131
rect 3467 4097 3476 4131
rect 3424 4088 3476 4097
rect 3700 4131 3752 4140
rect 3700 4097 3709 4131
rect 3709 4097 3743 4131
rect 3743 4097 3752 4131
rect 3700 4088 3752 4097
rect 4160 4020 4212 4072
rect 6368 4088 6420 4140
rect 6552 4131 6604 4140
rect 6552 4097 6561 4131
rect 6561 4097 6595 4131
rect 6595 4097 6604 4131
rect 6552 4088 6604 4097
rect 7288 4088 7340 4140
rect 7564 4088 7616 4140
rect 7748 4088 7800 4140
rect 7840 4088 7892 4140
rect 11244 4156 11296 4208
rect 13728 4156 13780 4208
rect 14832 4156 14884 4208
rect 21364 4156 21416 4208
rect 8576 4088 8628 4140
rect 13820 4088 13872 4140
rect 6460 4020 6512 4072
rect 3516 3884 3568 3936
rect 3608 3927 3660 3936
rect 3608 3893 3617 3927
rect 3617 3893 3651 3927
rect 3651 3893 3660 3927
rect 3608 3884 3660 3893
rect 3884 3927 3936 3936
rect 3884 3893 3893 3927
rect 3893 3893 3927 3927
rect 3927 3893 3936 3927
rect 3884 3884 3936 3893
rect 4436 3927 4488 3936
rect 4436 3893 4445 3927
rect 4445 3893 4479 3927
rect 4479 3893 4488 3927
rect 4436 3884 4488 3893
rect 14372 4020 14424 4072
rect 9680 3952 9732 4004
rect 14556 4088 14608 4140
rect 15844 4088 15896 4140
rect 22836 4088 22888 4140
rect 27344 4088 27396 4140
rect 5632 3884 5684 3936
rect 7196 3884 7248 3936
rect 7472 3884 7524 3936
rect 7656 3884 7708 3936
rect 8024 3884 8076 3936
rect 13636 3884 13688 3936
rect 21824 4020 21876 4072
rect 23940 4020 23992 4072
rect 27896 4020 27948 4072
rect 22284 3952 22336 4004
rect 24676 3952 24728 4004
rect 29552 4131 29604 4140
rect 29552 4097 29561 4131
rect 29561 4097 29595 4131
rect 29595 4097 29604 4131
rect 29552 4088 29604 4097
rect 30564 4088 30616 4140
rect 28448 4063 28500 4072
rect 28448 4029 28457 4063
rect 28457 4029 28491 4063
rect 28491 4029 28500 4063
rect 28448 4020 28500 4029
rect 28908 4020 28960 4072
rect 28724 3952 28776 4004
rect 32864 3995 32916 4004
rect 32864 3961 32873 3995
rect 32873 3961 32907 3995
rect 32907 3961 32916 3995
rect 32864 3952 32916 3961
rect 14648 3927 14700 3936
rect 14648 3893 14657 3927
rect 14657 3893 14691 3927
rect 14691 3893 14700 3927
rect 14648 3884 14700 3893
rect 15660 3884 15712 3936
rect 25504 3884 25556 3936
rect 27528 3927 27580 3936
rect 27528 3893 27537 3927
rect 27537 3893 27571 3927
rect 27571 3893 27580 3927
rect 27528 3884 27580 3893
rect 27712 3884 27764 3936
rect 27896 3884 27948 3936
rect 28816 3884 28868 3936
rect 29184 3927 29236 3936
rect 29184 3893 29193 3927
rect 29193 3893 29227 3927
rect 29227 3893 29236 3927
rect 29184 3884 29236 3893
rect 32496 3927 32548 3936
rect 32496 3893 32505 3927
rect 32505 3893 32539 3927
rect 32539 3893 32548 3927
rect 32496 3884 32548 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 13950 3782 14002 3834
rect 14014 3782 14066 3834
rect 14078 3782 14130 3834
rect 14142 3782 14194 3834
rect 14206 3782 14258 3834
rect 19950 3782 20002 3834
rect 20014 3782 20066 3834
rect 20078 3782 20130 3834
rect 20142 3782 20194 3834
rect 20206 3782 20258 3834
rect 25950 3782 26002 3834
rect 26014 3782 26066 3834
rect 26078 3782 26130 3834
rect 26142 3782 26194 3834
rect 26206 3782 26258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 3700 3680 3752 3732
rect 6736 3680 6788 3732
rect 7656 3680 7708 3732
rect 18972 3680 19024 3732
rect 3424 3612 3476 3664
rect 6920 3612 6972 3664
rect 7012 3612 7064 3664
rect 16580 3612 16632 3664
rect 17132 3612 17184 3664
rect 24124 3723 24176 3732
rect 24124 3689 24133 3723
rect 24133 3689 24167 3723
rect 24167 3689 24176 3723
rect 24124 3680 24176 3689
rect 26056 3680 26108 3732
rect 26884 3680 26936 3732
rect 28908 3680 28960 3732
rect 20904 3612 20956 3664
rect 2872 3544 2924 3596
rect 7288 3544 7340 3596
rect 7380 3544 7432 3596
rect 8392 3544 8444 3596
rect 13728 3544 13780 3596
rect 19708 3544 19760 3596
rect 20720 3587 20772 3596
rect 20720 3553 20729 3587
rect 20729 3553 20763 3587
rect 20763 3553 20772 3587
rect 24768 3612 24820 3664
rect 20720 3544 20772 3553
rect 7104 3476 7156 3528
rect 8760 3476 8812 3528
rect 13636 3476 13688 3528
rect 17776 3476 17828 3528
rect 22376 3544 22428 3596
rect 23388 3544 23440 3596
rect 2596 3408 2648 3460
rect 4896 3408 4948 3460
rect 6552 3408 6604 3460
rect 9404 3408 9456 3460
rect 14372 3408 14424 3460
rect 17408 3408 17460 3460
rect 17500 3408 17552 3460
rect 20352 3408 20404 3460
rect 2504 3383 2556 3392
rect 2504 3349 2513 3383
rect 2513 3349 2547 3383
rect 2547 3349 2556 3383
rect 2504 3340 2556 3349
rect 7380 3383 7432 3392
rect 7380 3349 7389 3383
rect 7389 3349 7423 3383
rect 7423 3349 7432 3383
rect 7380 3340 7432 3349
rect 12716 3340 12768 3392
rect 17592 3340 17644 3392
rect 17684 3340 17736 3392
rect 19156 3340 19208 3392
rect 19616 3340 19668 3392
rect 21916 3476 21968 3528
rect 25320 3544 25372 3596
rect 26148 3544 26200 3596
rect 26792 3544 26844 3596
rect 21640 3340 21692 3392
rect 22100 3340 22152 3392
rect 22192 3383 22244 3392
rect 22192 3349 22201 3383
rect 22201 3349 22235 3383
rect 22235 3349 22244 3383
rect 22192 3340 22244 3349
rect 23572 3383 23624 3392
rect 23572 3349 23581 3383
rect 23581 3349 23615 3383
rect 23615 3349 23624 3383
rect 23572 3340 23624 3349
rect 24860 3476 24912 3528
rect 26332 3476 26384 3528
rect 26516 3476 26568 3528
rect 26884 3519 26936 3528
rect 26884 3485 26893 3519
rect 26893 3485 26927 3519
rect 26927 3485 26936 3519
rect 26884 3476 26936 3485
rect 27436 3519 27488 3528
rect 27436 3485 27445 3519
rect 27445 3485 27479 3519
rect 27479 3485 27488 3519
rect 27436 3476 27488 3485
rect 24584 3383 24636 3392
rect 24584 3349 24593 3383
rect 24593 3349 24627 3383
rect 24627 3349 24636 3383
rect 24584 3340 24636 3349
rect 25044 3408 25096 3460
rect 25320 3340 25372 3392
rect 25780 3340 25832 3392
rect 26700 3383 26752 3392
rect 26700 3349 26709 3383
rect 26709 3349 26743 3383
rect 26743 3349 26752 3383
rect 26700 3340 26752 3349
rect 26792 3340 26844 3392
rect 27804 3544 27856 3596
rect 27896 3476 27948 3528
rect 28356 3476 28408 3528
rect 32864 3655 32916 3664
rect 32864 3621 32873 3655
rect 32873 3621 32907 3655
rect 32907 3621 32916 3655
rect 32864 3612 32916 3621
rect 30380 3544 30432 3596
rect 28172 3340 28224 3392
rect 28540 3383 28592 3392
rect 28540 3349 28549 3383
rect 28549 3349 28583 3383
rect 28583 3349 28592 3383
rect 28540 3340 28592 3349
rect 33416 3340 33468 3392
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 9010 3238 9062 3290
rect 9074 3238 9126 3290
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 15010 3238 15062 3290
rect 15074 3238 15126 3290
rect 15138 3238 15190 3290
rect 15202 3238 15254 3290
rect 15266 3238 15318 3290
rect 21010 3238 21062 3290
rect 21074 3238 21126 3290
rect 21138 3238 21190 3290
rect 21202 3238 21254 3290
rect 21266 3238 21318 3290
rect 27010 3238 27062 3290
rect 27074 3238 27126 3290
rect 27138 3238 27190 3290
rect 27202 3238 27254 3290
rect 27266 3238 27318 3290
rect 33010 3238 33062 3290
rect 33074 3238 33126 3290
rect 33138 3238 33190 3290
rect 33202 3238 33254 3290
rect 33266 3238 33318 3290
rect 2412 3136 2464 3188
rect 4528 3136 4580 3188
rect 10140 3136 10192 3188
rect 15936 3136 15988 3188
rect 17592 3136 17644 3188
rect 11796 3068 11848 3120
rect 15476 3043 15528 3052
rect 15476 3009 15485 3043
rect 15485 3009 15519 3043
rect 15519 3009 15528 3043
rect 15476 3000 15528 3009
rect 3884 2932 3936 2984
rect 16028 3000 16080 3052
rect 16764 3043 16816 3052
rect 16764 3009 16773 3043
rect 16773 3009 16807 3043
rect 16807 3009 16816 3043
rect 16764 3000 16816 3009
rect 2688 2864 2740 2916
rect 14832 2864 14884 2916
rect 15936 2932 15988 2984
rect 17408 3000 17460 3052
rect 18972 3043 19024 3052
rect 18972 3009 18981 3043
rect 18981 3009 19015 3043
rect 19015 3009 19024 3043
rect 18972 3000 19024 3009
rect 19248 3000 19300 3052
rect 19708 3043 19760 3052
rect 19708 3009 19717 3043
rect 19717 3009 19751 3043
rect 19751 3009 19760 3043
rect 19708 3000 19760 3009
rect 20444 3043 20496 3052
rect 20444 3009 20453 3043
rect 20453 3009 20487 3043
rect 20487 3009 20496 3043
rect 20444 3000 20496 3009
rect 22008 3136 22060 3188
rect 23664 3136 23716 3188
rect 24768 3136 24820 3188
rect 27068 3136 27120 3188
rect 27528 3136 27580 3188
rect 27804 3136 27856 3188
rect 32864 3179 32916 3188
rect 32864 3145 32873 3179
rect 32873 3145 32907 3179
rect 32907 3145 32916 3179
rect 32864 3136 32916 3145
rect 17224 2932 17276 2984
rect 20352 2932 20404 2984
rect 20628 2932 20680 2984
rect 21824 3043 21876 3052
rect 21824 3009 21833 3043
rect 21833 3009 21867 3043
rect 21867 3009 21876 3043
rect 21824 3000 21876 3009
rect 22284 3000 22336 3052
rect 22836 3043 22888 3052
rect 22836 3009 22845 3043
rect 22845 3009 22879 3043
rect 22879 3009 22888 3043
rect 22836 3000 22888 3009
rect 23204 3043 23256 3052
rect 23204 3009 23213 3043
rect 23213 3009 23247 3043
rect 23247 3009 23256 3043
rect 23204 3000 23256 3009
rect 22928 2932 22980 2984
rect 23940 3043 23992 3052
rect 23940 3009 23949 3043
rect 23949 3009 23983 3043
rect 23983 3009 23992 3043
rect 23940 3000 23992 3009
rect 24676 3043 24728 3052
rect 24676 3009 24685 3043
rect 24685 3009 24719 3043
rect 24719 3009 24728 3043
rect 24676 3000 24728 3009
rect 25044 3043 25096 3052
rect 25044 3009 25053 3043
rect 25053 3009 25087 3043
rect 25087 3009 25096 3043
rect 25044 3000 25096 3009
rect 25504 3000 25556 3052
rect 25780 3043 25832 3052
rect 25780 3009 25789 3043
rect 25789 3009 25823 3043
rect 25823 3009 25832 3043
rect 25780 3000 25832 3009
rect 28448 3068 28500 3120
rect 27804 3043 27856 3052
rect 27804 3009 27813 3043
rect 27813 3009 27847 3043
rect 27847 3009 27856 3043
rect 27804 3000 27856 3009
rect 31668 3043 31720 3052
rect 31668 3009 31677 3043
rect 31677 3009 31711 3043
rect 31711 3009 31720 3043
rect 31668 3000 31720 3009
rect 16580 2864 16632 2916
rect 17776 2864 17828 2916
rect 17868 2864 17920 2916
rect 19064 2864 19116 2916
rect 19340 2864 19392 2916
rect 19708 2864 19760 2916
rect 19800 2864 19852 2916
rect 20536 2864 20588 2916
rect 21640 2864 21692 2916
rect 22468 2864 22520 2916
rect 23296 2864 23348 2916
rect 10600 2796 10652 2848
rect 12532 2796 12584 2848
rect 15384 2796 15436 2848
rect 15752 2796 15804 2848
rect 16120 2796 16172 2848
rect 16672 2796 16724 2848
rect 17040 2796 17092 2848
rect 17408 2796 17460 2848
rect 18880 2796 18932 2848
rect 19248 2796 19300 2848
rect 19616 2796 19668 2848
rect 20352 2796 20404 2848
rect 20720 2796 20772 2848
rect 21456 2796 21508 2848
rect 22744 2796 22796 2848
rect 24032 2864 24084 2916
rect 24400 2796 24452 2848
rect 28264 2864 28316 2916
rect 25780 2796 25832 2848
rect 28816 2796 28868 2848
rect 32404 2796 32456 2848
rect 32496 2839 32548 2848
rect 32496 2805 32505 2839
rect 32505 2805 32539 2839
rect 32539 2805 32548 2839
rect 32496 2796 32548 2805
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 13950 2694 14002 2746
rect 14014 2694 14066 2746
rect 14078 2694 14130 2746
rect 14142 2694 14194 2746
rect 14206 2694 14258 2746
rect 19950 2694 20002 2746
rect 20014 2694 20066 2746
rect 20078 2694 20130 2746
rect 20142 2694 20194 2746
rect 20206 2694 20258 2746
rect 25950 2694 26002 2746
rect 26014 2694 26066 2746
rect 26078 2694 26130 2746
rect 26142 2694 26194 2746
rect 26206 2694 26258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 3608 2592 3660 2644
rect 11060 2592 11112 2644
rect 2780 2524 2832 2576
rect 15476 2592 15528 2644
rect 18512 2592 18564 2644
rect 20168 2592 20220 2644
rect 21824 2592 21876 2644
rect 15568 2524 15620 2576
rect 16488 2524 16540 2576
rect 18144 2524 18196 2576
rect 19892 2524 19944 2576
rect 20904 2524 20956 2576
rect 3516 2456 3568 2508
rect 10416 2388 10468 2440
rect 13360 2388 13412 2440
rect 13452 2388 13504 2440
rect 4160 2320 4212 2372
rect 15476 2431 15528 2440
rect 15476 2397 15485 2431
rect 15485 2397 15519 2431
rect 15519 2397 15528 2431
rect 15476 2388 15528 2397
rect 16304 2456 16356 2508
rect 16212 2431 16264 2440
rect 16212 2397 16221 2431
rect 16221 2397 16255 2431
rect 16255 2397 16264 2431
rect 16212 2388 16264 2397
rect 16948 2431 17000 2440
rect 16948 2397 16957 2431
rect 16957 2397 16991 2431
rect 16991 2397 17000 2431
rect 16948 2388 17000 2397
rect 17316 2431 17368 2440
rect 17316 2397 17325 2431
rect 17325 2397 17359 2431
rect 17359 2397 17368 2431
rect 17316 2388 17368 2397
rect 17776 2456 17828 2508
rect 18052 2431 18104 2440
rect 18052 2397 18061 2431
rect 18061 2397 18095 2431
rect 18095 2397 18104 2431
rect 18052 2388 18104 2397
rect 18420 2431 18472 2440
rect 18420 2397 18429 2431
rect 18429 2397 18463 2431
rect 18463 2397 18472 2431
rect 18420 2388 18472 2397
rect 19064 2456 19116 2508
rect 19432 2456 19484 2508
rect 19340 2388 19392 2440
rect 19984 2431 20036 2440
rect 19984 2397 19993 2431
rect 19993 2397 20027 2431
rect 20027 2397 20036 2431
rect 19984 2388 20036 2397
rect 21272 2456 21324 2508
rect 22652 2592 22704 2644
rect 24216 2592 24268 2644
rect 25872 2592 25924 2644
rect 22192 2524 22244 2576
rect 23480 2524 23532 2576
rect 20812 2388 20864 2440
rect 10232 2252 10284 2304
rect 13084 2252 13136 2304
rect 15936 2320 15988 2372
rect 19064 2320 19116 2372
rect 16304 2252 16356 2304
rect 16856 2252 16908 2304
rect 17224 2252 17276 2304
rect 17592 2252 17644 2304
rect 17776 2252 17828 2304
rect 17960 2252 18012 2304
rect 18328 2252 18380 2304
rect 18696 2252 18748 2304
rect 20444 2320 20496 2372
rect 21732 2388 21784 2440
rect 22560 2431 22612 2440
rect 22560 2397 22569 2431
rect 22569 2397 22603 2431
rect 22603 2397 22612 2431
rect 22560 2388 22612 2397
rect 21456 2320 21508 2372
rect 20260 2252 20312 2304
rect 20996 2252 21048 2304
rect 21548 2252 21600 2304
rect 21732 2252 21784 2304
rect 23020 2388 23072 2440
rect 23572 2431 23624 2440
rect 23572 2397 23581 2431
rect 23581 2397 23615 2431
rect 23615 2397 23624 2431
rect 23572 2388 23624 2397
rect 23940 2431 23992 2440
rect 23940 2397 23949 2431
rect 23949 2397 23983 2431
rect 23983 2397 23992 2431
rect 23940 2388 23992 2397
rect 24492 2388 24544 2440
rect 23848 2320 23900 2372
rect 25320 2388 25372 2440
rect 27804 2524 27856 2576
rect 26792 2456 26844 2508
rect 26700 2388 26752 2440
rect 30932 2431 30984 2440
rect 30932 2397 30941 2431
rect 30941 2397 30975 2431
rect 30975 2397 30984 2431
rect 30932 2388 30984 2397
rect 31300 2431 31352 2440
rect 31300 2397 31309 2431
rect 31309 2397 31343 2431
rect 31343 2397 31352 2431
rect 31300 2388 31352 2397
rect 31668 2431 31720 2440
rect 31668 2397 31677 2431
rect 31677 2397 31711 2431
rect 31711 2397 31720 2431
rect 31668 2388 31720 2397
rect 32312 2431 32364 2440
rect 32312 2397 32321 2431
rect 32321 2397 32355 2431
rect 32355 2397 32364 2431
rect 32312 2388 32364 2397
rect 32864 2567 32916 2576
rect 32864 2533 32873 2567
rect 32873 2533 32907 2567
rect 32907 2533 32916 2567
rect 32864 2524 32916 2533
rect 23204 2252 23256 2304
rect 24584 2252 24636 2304
rect 31116 2295 31168 2304
rect 31116 2261 31125 2295
rect 31125 2261 31159 2295
rect 31159 2261 31168 2295
rect 31116 2252 31168 2261
rect 31484 2295 31536 2304
rect 31484 2261 31493 2295
rect 31493 2261 31527 2295
rect 31527 2261 31536 2295
rect 31484 2252 31536 2261
rect 31852 2295 31904 2304
rect 31852 2261 31861 2295
rect 31861 2261 31895 2295
rect 31895 2261 31904 2295
rect 31852 2252 31904 2261
rect 33416 2252 33468 2304
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 9010 2150 9062 2202
rect 9074 2150 9126 2202
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 15010 2150 15062 2202
rect 15074 2150 15126 2202
rect 15138 2150 15190 2202
rect 15202 2150 15254 2202
rect 15266 2150 15318 2202
rect 21010 2150 21062 2202
rect 21074 2150 21126 2202
rect 21138 2150 21190 2202
rect 21202 2150 21254 2202
rect 21266 2150 21318 2202
rect 27010 2150 27062 2202
rect 27074 2150 27126 2202
rect 27138 2150 27190 2202
rect 27202 2150 27254 2202
rect 27266 2150 27318 2202
rect 33010 2150 33062 2202
rect 33074 2150 33126 2202
rect 33138 2150 33190 2202
rect 33202 2150 33254 2202
rect 33266 2150 33318 2202
rect 11060 2048 11112 2100
rect 16212 2048 16264 2100
rect 16396 2048 16448 2100
rect 19984 2048 20036 2100
rect 22376 2048 22428 2100
rect 7472 1980 7524 2032
rect 18420 1980 18472 2032
rect 18604 1980 18656 2032
rect 22560 1980 22612 2032
rect 23572 2048 23624 2100
rect 28172 2048 28224 2100
rect 31300 1980 31352 2032
rect 17132 1912 17184 1964
rect 20444 1912 20496 1964
rect 22100 1912 22152 1964
rect 30932 1912 30984 1964
rect 7196 1844 7248 1896
rect 17316 1844 17368 1896
rect 19156 1844 19208 1896
rect 31668 1844 31720 1896
rect 8300 1776 8352 1828
rect 19340 1776 19392 1828
rect 24308 1776 24360 1828
rect 27712 1776 27764 1828
rect 7380 1708 7432 1760
rect 18052 1708 18104 1760
rect 4436 1640 4488 1692
rect 16948 1640 17000 1692
rect 14464 1572 14516 1624
rect 29184 1640 29236 1692
rect 27344 1572 27396 1624
rect 29644 1572 29696 1624
rect 15660 1504 15712 1556
rect 23020 1504 23072 1556
rect 28448 1504 28500 1556
rect 30840 1504 30892 1556
rect 14648 1436 14700 1488
rect 18604 1436 18656 1488
rect 19524 1436 19576 1488
rect 19892 1436 19944 1488
rect 21548 1436 21600 1488
rect 32312 1436 32364 1488
rect 19708 1368 19760 1420
rect 20260 1368 20312 1420
rect 21088 1368 21140 1420
rect 21732 1368 21784 1420
rect 27160 1368 27212 1420
rect 27620 1368 27672 1420
rect 28264 1368 28316 1420
rect 29920 1368 29972 1420
rect 9312 1300 9364 1352
rect 14556 1300 14608 1352
rect 9496 1232 9548 1284
rect 15844 1232 15896 1284
rect 14924 688 14976 740
rect 25504 688 25556 740
rect 14832 484 14884 536
rect 28540 484 28592 536
rect 14372 416 14424 468
rect 28356 416 28408 468
rect 12256 348 12308 400
rect 26516 348 26568 400
rect 13176 280 13228 332
rect 28724 280 28776 332
rect 12624 212 12676 264
rect 12808 144 12860 196
rect 15016 212 15068 264
rect 29552 212 29604 264
rect 13084 76 13136 128
rect 27252 144 27304 196
rect 27436 76 27488 128
rect 27804 76 27856 128
<< metal2 >>
rect 1490 11096 1546 11152
rect 2884 11110 3004 11138
rect 1306 9616 1362 9625
rect 1306 9551 1362 9560
rect 1124 7948 1176 7954
rect 1124 7890 1176 7896
rect 848 6996 900 7002
rect 848 6938 900 6944
rect 860 4729 888 6938
rect 846 4720 902 4729
rect 846 4655 902 4664
rect 1136 4185 1164 7890
rect 1216 7336 1268 7342
rect 1216 7278 1268 7284
rect 1228 4457 1256 7278
rect 1320 6798 1348 9551
rect 1504 8634 1532 11096
rect 2778 8800 2834 8809
rect 2778 8735 2834 8744
rect 1492 8628 1544 8634
rect 1492 8570 1544 8576
rect 2792 8401 2820 8735
rect 2884 8634 2912 11110
rect 2976 11098 3004 11110
rect 3054 11098 3110 11152
rect 2976 11096 3110 11098
rect 4618 11096 4674 11152
rect 6182 11096 6238 11152
rect 7746 11096 7802 11152
rect 9310 11096 9366 11152
rect 10874 11096 10930 11152
rect 12438 11096 12494 11152
rect 14002 11096 14058 11152
rect 15566 11096 15622 11152
rect 17130 11096 17186 11152
rect 18694 11096 18750 11152
rect 20258 11096 20314 11152
rect 21822 11096 21878 11152
rect 23386 11096 23442 11152
rect 24950 11096 25006 11152
rect 26514 11096 26570 11152
rect 28078 11096 28134 11152
rect 29642 11096 29698 11152
rect 31206 11096 31262 11152
rect 32770 11096 32826 11152
rect 2976 11070 3096 11096
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 4632 8634 4660 11096
rect 6196 8634 6224 11096
rect 7760 8634 7788 11096
rect 9324 8922 9352 11096
rect 9324 8894 9444 8922
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 8036 8498 8064 8774
rect 9010 8732 9318 8741
rect 9010 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9176 8732
rect 9232 8730 9256 8732
rect 9312 8730 9318 8732
rect 9072 8678 9074 8730
rect 9254 8678 9256 8730
rect 9010 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9176 8678
rect 9232 8676 9256 8678
rect 9312 8676 9318 8678
rect 9010 8667 9318 8676
rect 9416 8634 9444 8894
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 2778 8392 2834 8401
rect 10888 8362 10916 11096
rect 11244 8900 11296 8906
rect 11244 8842 11296 8848
rect 11060 8560 11112 8566
rect 11060 8502 11112 8508
rect 2778 8327 2834 8336
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 5540 8288 5592 8294
rect 1766 8256 1822 8265
rect 5540 8230 5592 8236
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 1766 8191 1822 8200
rect 1400 7744 1452 7750
rect 1400 7686 1452 7692
rect 1308 6792 1360 6798
rect 1308 6734 1360 6740
rect 1412 5658 1440 7686
rect 1676 7268 1728 7274
rect 1676 7210 1728 7216
rect 1320 5630 1440 5658
rect 1320 5001 1348 5630
rect 1306 4992 1362 5001
rect 1306 4927 1362 4936
rect 1306 4584 1362 4593
rect 1306 4519 1362 4528
rect 1214 4448 1270 4457
rect 1214 4383 1270 4392
rect 1122 4176 1178 4185
rect 1122 4111 1178 4120
rect 1320 2825 1348 4519
rect 1688 3913 1716 7210
rect 1780 6866 1808 8191
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 2594 7984 2650 7993
rect 2594 7919 2650 7928
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 2608 6458 2636 7919
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 5552 7546 5580 8230
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 9010 7644 9318 7653
rect 9010 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9176 7644
rect 9232 7642 9256 7644
rect 9312 7642 9318 7644
rect 9072 7590 9074 7642
rect 9254 7590 9256 7642
rect 9010 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9176 7590
rect 9232 7588 9256 7590
rect 9312 7588 9318 7590
rect 9010 7579 9318 7588
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 9508 7206 9536 8230
rect 11072 7546 11100 8502
rect 11256 8498 11284 8842
rect 12452 8634 12480 11096
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12820 8498 12848 8978
rect 14016 8634 14044 11096
rect 14372 9104 14424 9110
rect 14372 9046 14424 9052
rect 14738 9072 14794 9081
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 14384 8498 14412 9046
rect 14738 9007 14794 9016
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 12360 7410 12388 7686
rect 13832 7546 13860 8298
rect 13950 8188 14258 8197
rect 13950 8186 13956 8188
rect 14012 8186 14036 8188
rect 14092 8186 14116 8188
rect 14172 8186 14196 8188
rect 14252 8186 14258 8188
rect 14012 8134 14014 8186
rect 14194 8134 14196 8186
rect 13950 8132 13956 8134
rect 14012 8132 14036 8134
rect 14092 8132 14116 8134
rect 14172 8132 14196 8134
rect 14252 8132 14258 8134
rect 13950 8123 14258 8132
rect 14372 7880 14424 7886
rect 14372 7822 14424 7828
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 14384 7410 14412 7822
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 2688 6928 2740 6934
rect 2688 6870 2740 6876
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 1766 6080 1822 6089
rect 1766 6015 1822 6024
rect 1780 5681 1808 6015
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 1766 5672 1822 5681
rect 1766 5607 1822 5616
rect 2700 5273 2728 6870
rect 2870 6624 2926 6633
rect 2870 6559 2926 6568
rect 2780 6248 2832 6254
rect 2884 6225 2912 6559
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 9010 6556 9318 6565
rect 9010 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9176 6556
rect 9232 6554 9256 6556
rect 9312 6554 9318 6556
rect 9072 6502 9074 6554
rect 9254 6502 9256 6554
rect 9010 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9176 6502
rect 9232 6500 9256 6502
rect 9312 6500 9318 6502
rect 9010 6491 9318 6500
rect 2780 6190 2832 6196
rect 2870 6216 2926 6225
rect 2792 5545 2820 6190
rect 2870 6151 2926 6160
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 9600 5846 9628 7346
rect 13950 7100 14258 7109
rect 13950 7098 13956 7100
rect 14012 7098 14036 7100
rect 14092 7098 14116 7100
rect 14172 7098 14196 7100
rect 14252 7098 14258 7100
rect 14012 7046 14014 7098
rect 14194 7046 14196 7098
rect 13950 7044 13956 7046
rect 14012 7044 14036 7046
rect 14092 7044 14116 7046
rect 14172 7044 14196 7046
rect 14252 7044 14258 7046
rect 13950 7035 14258 7044
rect 13950 6012 14258 6021
rect 13950 6010 13956 6012
rect 14012 6010 14036 6012
rect 14092 6010 14116 6012
rect 14172 6010 14196 6012
rect 14252 6010 14258 6012
rect 14012 5958 14014 6010
rect 14194 5958 14196 6010
rect 13950 5956 13956 5958
rect 14012 5956 14036 5958
rect 14092 5956 14116 5958
rect 14172 5956 14196 5958
rect 14252 5956 14258 5958
rect 13950 5947 14258 5956
rect 9588 5840 9640 5846
rect 9588 5782 9640 5788
rect 2778 5536 2834 5545
rect 2778 5471 2834 5480
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 9010 5468 9318 5477
rect 9010 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9176 5468
rect 9232 5466 9256 5468
rect 9312 5466 9318 5468
rect 9072 5414 9074 5466
rect 9254 5414 9256 5466
rect 9010 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9176 5414
rect 9232 5412 9256 5414
rect 9312 5412 9318 5414
rect 9010 5403 9318 5412
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 3424 5296 3476 5302
rect 2686 5264 2742 5273
rect 3424 5238 3476 5244
rect 7380 5296 7432 5302
rect 7380 5238 7432 5244
rect 2686 5199 2742 5208
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 3160 4826 3188 5170
rect 3436 4826 3464 5238
rect 7392 4826 7420 5238
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3424 4820 3476 4826
rect 3424 4762 3476 4768
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 2688 4276 2740 4282
rect 2688 4218 2740 4224
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 1674 3904 1730 3913
rect 1674 3839 1730 3848
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 2424 3194 2452 4082
rect 2502 3496 2558 3505
rect 2608 3466 2636 4082
rect 2502 3431 2558 3440
rect 2596 3460 2648 3466
rect 2516 3398 2544 3431
rect 2596 3402 2648 3408
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 2700 2922 2728 4218
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 2780 4004 2832 4010
rect 2780 3946 2832 3952
rect 2688 2916 2740 2922
rect 2688 2858 2740 2864
rect 1306 2816 1362 2825
rect 1306 2751 1362 2760
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 2792 2582 2820 3946
rect 2884 3602 2912 4014
rect 3436 3670 3464 4082
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3608 3936 3660 3942
rect 3608 3878 3660 3884
rect 3424 3664 3476 3670
rect 3424 3606 3476 3612
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 2870 3360 2926 3369
rect 2870 3295 2926 3304
rect 2884 2961 2912 3295
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 2870 2952 2926 2961
rect 2870 2887 2926 2896
rect 2780 2576 2832 2582
rect 2780 2518 2832 2524
rect 3528 2514 3556 3878
rect 3620 2650 3648 3878
rect 3712 3738 3740 4082
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3700 3732 3752 3738
rect 3700 3674 3752 3680
rect 3896 2990 3924 3878
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 3608 2644 3660 2650
rect 3608 2586 3660 2592
rect 3516 2508 3568 2514
rect 3516 2450 3568 2456
rect 4172 2378 4200 4014
rect 4436 3936 4488 3942
rect 4436 3878 4488 3884
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 2870 2272 2926 2281
rect 2870 2207 2926 2216
rect 2884 1873 2912 2207
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 2870 1864 2926 1873
rect 2870 1799 2926 1808
rect 4448 1698 4476 3878
rect 4896 3460 4948 3466
rect 4896 3402 4948 3408
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4436 1692 4488 1698
rect 4436 1634 4488 1640
rect 4540 1329 4568 3130
rect 4526 1320 4582 1329
rect 4526 1255 4582 1264
rect 4908 105 4936 3402
rect 4894 96 4950 105
rect 5644 56 5672 3878
rect 5828 56 5856 4558
rect 6000 4548 6052 4554
rect 6000 4490 6052 4496
rect 6012 56 6040 4490
rect 6196 56 6224 4626
rect 8852 4616 8904 4622
rect 8852 4558 8904 4564
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6380 56 6408 4082
rect 6460 4072 6512 4078
rect 6460 4014 6512 4020
rect 6472 82 6500 4014
rect 6564 3466 6592 4082
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6552 3460 6604 3466
rect 6552 3402 6604 3408
rect 6472 56 6592 82
rect 6748 56 6776 3674
rect 7024 3670 7052 4218
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 7012 3664 7064 3670
rect 7012 3606 7064 3612
rect 6932 56 6960 3606
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 7116 56 7144 3470
rect 7208 1902 7236 3878
rect 7300 3720 7328 4082
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7300 3692 7420 3720
rect 7392 3602 7420 3692
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7196 1896 7248 1902
rect 7196 1838 7248 1844
rect 7300 56 7328 3538
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7392 1766 7420 3334
rect 7484 2038 7512 3878
rect 7472 2032 7524 2038
rect 7472 1974 7524 1980
rect 7380 1760 7432 1766
rect 7380 1702 7432 1708
rect 7470 1320 7526 1329
rect 7470 1255 7526 1264
rect 7484 56 7512 1255
rect 7576 218 7604 4082
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7668 3738 7696 3878
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 7760 1986 7788 4082
rect 7852 2122 7880 4082
rect 8036 3998 8340 4026
rect 8036 3942 8064 3998
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 8312 3720 8340 3998
rect 8220 3692 8340 3720
rect 8220 2836 8248 3692
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 8220 2808 8340 2836
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 7852 2094 8248 2122
rect 7760 1958 8064 1986
rect 7576 190 7880 218
rect 7654 96 7710 105
rect 4894 31 4950 40
rect 5630 0 5686 56
rect 5814 0 5870 56
rect 5998 0 6054 56
rect 6182 0 6238 56
rect 6366 0 6422 56
rect 6472 54 6606 56
rect 6550 0 6606 54
rect 6734 0 6790 56
rect 6918 0 6974 56
rect 7102 0 7158 56
rect 7286 0 7342 56
rect 7470 0 7526 56
rect 7852 56 7880 190
rect 8036 56 8064 1958
rect 8220 56 8248 2094
rect 8312 1834 8340 2808
rect 8300 1828 8352 1834
rect 8300 1770 8352 1776
rect 8404 56 8432 3538
rect 8588 56 8616 4082
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8772 56 8800 3470
rect 8864 82 8892 4558
rect 9010 4380 9318 4389
rect 9010 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9176 4380
rect 9232 4378 9256 4380
rect 9312 4378 9318 4380
rect 9072 4326 9074 4378
rect 9254 4326 9256 4378
rect 9010 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9176 4326
rect 9232 4324 9256 4326
rect 9312 4324 9318 4326
rect 9010 4315 9318 4324
rect 9680 4004 9732 4010
rect 9680 3946 9732 3952
rect 9404 3460 9456 3466
rect 9404 3402 9456 3408
rect 9010 3292 9318 3301
rect 9010 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9176 3292
rect 9232 3290 9256 3292
rect 9312 3290 9318 3292
rect 9072 3238 9074 3290
rect 9254 3238 9256 3290
rect 9010 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9176 3238
rect 9232 3236 9256 3238
rect 9312 3236 9318 3238
rect 9010 3227 9318 3236
rect 9010 2204 9318 2213
rect 9010 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9176 2204
rect 9232 2202 9256 2204
rect 9312 2202 9318 2204
rect 9072 2150 9074 2202
rect 9254 2150 9256 2202
rect 9010 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9176 2150
rect 9232 2148 9256 2150
rect 9312 2148 9318 2150
rect 9010 2139 9318 2148
rect 9416 1714 9444 3402
rect 9140 1686 9444 1714
rect 8864 56 8984 82
rect 9140 56 9168 1686
rect 9312 1352 9364 1358
rect 9312 1294 9364 1300
rect 9324 56 9352 1294
rect 9496 1284 9548 1290
rect 9496 1226 9548 1232
rect 9508 56 9536 1226
rect 9692 56 9720 3946
rect 9862 2136 9918 2145
rect 9862 2071 9918 2080
rect 9876 56 9904 2071
rect 10060 56 10088 5170
rect 13268 5160 13320 5166
rect 11058 5128 11114 5137
rect 13268 5102 13320 5108
rect 11058 5063 11114 5072
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 10140 4480 10192 4486
rect 10140 4422 10192 4428
rect 10152 3194 10180 4422
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10600 2848 10652 2854
rect 10600 2790 10652 2796
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 10244 56 10272 2246
rect 10428 56 10456 2382
rect 10612 56 10640 2790
rect 10796 56 10824 4218
rect 10980 56 11008 4762
rect 11072 4486 11100 5063
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 12084 4826 12112 4966
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 13280 4758 13308 5102
rect 11704 4752 11756 4758
rect 11610 4720 11666 4729
rect 11520 4684 11572 4690
rect 11704 4694 11756 4700
rect 13268 4752 13320 4758
rect 13268 4694 13320 4700
rect 11610 4655 11666 4664
rect 11520 4626 11572 4632
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11072 2106 11100 2586
rect 11060 2100 11112 2106
rect 11060 2042 11112 2048
rect 11164 56 11192 4490
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 11256 4214 11284 4422
rect 11244 4208 11296 4214
rect 11244 4150 11296 4156
rect 11348 56 11376 4558
rect 11532 56 11560 4626
rect 11624 4486 11652 4655
rect 11612 4480 11664 4486
rect 11612 4422 11664 4428
rect 11716 56 11744 4694
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 11796 4480 11848 4486
rect 11796 4422 11848 4428
rect 11808 3126 11836 4422
rect 11796 3120 11848 3126
rect 11796 3062 11848 3068
rect 11992 82 12020 4626
rect 12256 4616 12308 4622
rect 12256 4558 12308 4564
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 12072 4548 12124 4554
rect 12072 4490 12124 4496
rect 11900 56 12020 82
rect 12084 56 12112 4490
rect 12268 4282 12296 4558
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12452 4282 12480 4422
rect 12256 4276 12308 4282
rect 12256 4218 12308 4224
rect 12440 4276 12492 4282
rect 12440 4218 12492 4224
rect 12544 2854 12572 4558
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 12728 3398 12756 4422
rect 12716 3392 12768 3398
rect 12716 3334 12768 3340
rect 12532 2848 12584 2854
rect 12532 2790 12584 2796
rect 12438 2408 12494 2417
rect 12438 2343 12494 2352
rect 12256 400 12308 406
rect 12256 342 12308 348
rect 12268 56 12296 342
rect 12452 56 12480 2343
rect 13096 2310 13124 4558
rect 13372 2446 13400 4558
rect 13464 2446 13492 5306
rect 14752 5234 14780 9007
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14844 7546 14872 8774
rect 15010 8732 15318 8741
rect 15010 8730 15016 8732
rect 15072 8730 15096 8732
rect 15152 8730 15176 8732
rect 15232 8730 15256 8732
rect 15312 8730 15318 8732
rect 15072 8678 15074 8730
rect 15254 8678 15256 8730
rect 15010 8676 15016 8678
rect 15072 8676 15096 8678
rect 15152 8676 15176 8678
rect 15232 8676 15256 8678
rect 15312 8676 15318 8678
rect 15010 8667 15318 8676
rect 15580 8634 15608 11096
rect 16946 9344 17002 9353
rect 16946 9279 17002 9288
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 16580 8016 16632 8022
rect 16580 7958 16632 7964
rect 15010 7644 15318 7653
rect 15010 7642 15016 7644
rect 15072 7642 15096 7644
rect 15152 7642 15176 7644
rect 15232 7642 15256 7644
rect 15312 7642 15318 7644
rect 15072 7590 15074 7642
rect 15254 7590 15256 7642
rect 15010 7588 15016 7590
rect 15072 7588 15096 7590
rect 15152 7588 15176 7590
rect 15232 7588 15256 7590
rect 15312 7588 15318 7590
rect 15010 7579 15318 7588
rect 14832 7540 14884 7546
rect 14832 7482 14884 7488
rect 15474 7440 15530 7449
rect 14924 7404 14976 7410
rect 15474 7375 15530 7384
rect 14924 7346 14976 7352
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 13648 4622 13676 5170
rect 13950 4924 14258 4933
rect 13950 4922 13956 4924
rect 14012 4922 14036 4924
rect 14092 4922 14116 4924
rect 14172 4922 14196 4924
rect 14252 4922 14258 4924
rect 14012 4870 14014 4922
rect 14194 4870 14196 4922
rect 13950 4868 13956 4870
rect 14012 4868 14036 4870
rect 14092 4868 14116 4870
rect 14172 4868 14196 4870
rect 14252 4868 14258 4870
rect 13950 4859 14258 4868
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14844 4214 14872 4422
rect 13728 4208 13780 4214
rect 13728 4150 13780 4156
rect 14832 4208 14884 4214
rect 14832 4150 14884 4156
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13648 3534 13676 3878
rect 13740 3602 13768 4150
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 13452 2440 13504 2446
rect 13452 2382 13504 2388
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 13832 2145 13860 4082
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 13950 3836 14258 3845
rect 13950 3834 13956 3836
rect 14012 3834 14036 3836
rect 14092 3834 14116 3836
rect 14172 3834 14196 3836
rect 14252 3834 14258 3836
rect 14012 3782 14014 3834
rect 14194 3782 14196 3834
rect 13950 3780 13956 3782
rect 14012 3780 14036 3782
rect 14092 3780 14116 3782
rect 14172 3780 14196 3782
rect 14252 3780 14258 3782
rect 13950 3771 14258 3780
rect 14384 3466 14412 4014
rect 14462 3904 14518 3913
rect 14462 3839 14518 3848
rect 14372 3460 14424 3466
rect 14372 3402 14424 3408
rect 14476 2774 14504 3839
rect 13950 2748 14258 2757
rect 13950 2746 13956 2748
rect 14012 2746 14036 2748
rect 14092 2746 14116 2748
rect 14172 2746 14196 2748
rect 14252 2746 14258 2748
rect 14012 2694 14014 2746
rect 14194 2694 14196 2746
rect 13950 2692 13956 2694
rect 14012 2692 14036 2694
rect 14092 2692 14116 2694
rect 14172 2692 14196 2694
rect 14252 2692 14258 2694
rect 13950 2683 14258 2692
rect 14292 2746 14504 2774
rect 13818 2136 13874 2145
rect 13818 2071 13874 2080
rect 13726 640 13782 649
rect 13726 575 13782 584
rect 13542 504 13598 513
rect 13542 439 13598 448
rect 13358 368 13414 377
rect 13176 332 13228 338
rect 13358 303 13414 312
rect 13176 274 13228 280
rect 12624 264 12676 270
rect 12624 206 12676 212
rect 12636 56 12664 206
rect 12808 196 12860 202
rect 12808 138 12860 144
rect 13004 190 13124 218
rect 12820 56 12848 138
rect 13004 56 13032 190
rect 13096 134 13124 190
rect 13084 128 13136 134
rect 13084 70 13136 76
rect 13188 56 13216 274
rect 13372 56 13400 303
rect 13556 56 13584 439
rect 13740 56 13768 575
rect 13910 232 13966 241
rect 14292 218 14320 2746
rect 14464 1624 14516 1630
rect 14464 1566 14516 1572
rect 14372 468 14424 474
rect 14372 410 14424 416
rect 13910 167 13966 176
rect 14200 190 14320 218
rect 13924 56 13952 167
rect 14200 82 14228 190
rect 14384 82 14412 410
rect 14108 56 14228 82
rect 14292 56 14412 82
rect 14476 56 14504 1566
rect 14568 1358 14596 4082
rect 14738 4040 14794 4049
rect 14738 3975 14794 3984
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14660 1494 14688 3878
rect 14648 1488 14700 1494
rect 14648 1430 14700 1436
rect 14556 1352 14608 1358
rect 14556 1294 14608 1300
rect 14752 82 14780 3975
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 14844 2825 14872 2858
rect 14830 2816 14886 2825
rect 14830 2751 14886 2760
rect 14936 746 14964 7346
rect 15010 6556 15318 6565
rect 15010 6554 15016 6556
rect 15072 6554 15096 6556
rect 15152 6554 15176 6556
rect 15232 6554 15256 6556
rect 15312 6554 15318 6556
rect 15072 6502 15074 6554
rect 15254 6502 15256 6554
rect 15010 6500 15016 6502
rect 15072 6500 15096 6502
rect 15152 6500 15176 6502
rect 15232 6500 15256 6502
rect 15312 6500 15318 6502
rect 15010 6491 15318 6500
rect 15108 6384 15160 6390
rect 15106 6352 15108 6361
rect 15160 6352 15162 6361
rect 15106 6287 15162 6296
rect 15010 5468 15318 5477
rect 15010 5466 15016 5468
rect 15072 5466 15096 5468
rect 15152 5466 15176 5468
rect 15232 5466 15256 5468
rect 15312 5466 15318 5468
rect 15072 5414 15074 5466
rect 15254 5414 15256 5466
rect 15010 5412 15016 5414
rect 15072 5412 15096 5414
rect 15152 5412 15176 5414
rect 15232 5412 15256 5414
rect 15312 5412 15318 5414
rect 15010 5403 15318 5412
rect 15200 5296 15252 5302
rect 15488 5250 15516 7375
rect 16486 7304 16542 7313
rect 16486 7239 16542 7248
rect 15750 6896 15806 6905
rect 16500 6866 16528 7239
rect 15750 6831 15806 6840
rect 16488 6860 16540 6866
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 15580 5370 15608 6394
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 15200 5238 15252 5244
rect 15212 4486 15240 5238
rect 15396 5222 15516 5250
rect 15660 5296 15712 5302
rect 15660 5238 15712 5244
rect 15396 4826 15424 5222
rect 15672 5137 15700 5238
rect 15658 5128 15714 5137
rect 15476 5092 15528 5098
rect 15658 5063 15714 5072
rect 15476 5034 15528 5040
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 15010 4380 15318 4389
rect 15010 4378 15016 4380
rect 15072 4378 15096 4380
rect 15152 4378 15176 4380
rect 15232 4378 15256 4380
rect 15312 4378 15318 4380
rect 15072 4326 15074 4378
rect 15254 4326 15256 4378
rect 15010 4324 15016 4326
rect 15072 4324 15096 4326
rect 15152 4324 15176 4326
rect 15232 4324 15256 4326
rect 15312 4324 15318 4326
rect 15010 4315 15318 4324
rect 15010 3292 15318 3301
rect 15010 3290 15016 3292
rect 15072 3290 15096 3292
rect 15152 3290 15176 3292
rect 15232 3290 15256 3292
rect 15312 3290 15318 3292
rect 15072 3238 15074 3290
rect 15254 3238 15256 3290
rect 15010 3236 15016 3238
rect 15072 3236 15096 3238
rect 15152 3236 15176 3238
rect 15232 3236 15256 3238
rect 15312 3236 15318 3238
rect 15010 3227 15318 3236
rect 15488 3058 15516 5034
rect 15764 4622 15792 6831
rect 16488 6802 16540 6808
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 16132 6254 16160 6598
rect 16120 6248 16172 6254
rect 16120 6190 16172 6196
rect 16210 6216 16266 6225
rect 16210 6151 16266 6160
rect 15934 5264 15990 5273
rect 15934 5199 15990 5208
rect 15948 4826 15976 5199
rect 16224 4826 16252 6151
rect 16394 5672 16450 5681
rect 16592 5658 16620 7958
rect 16394 5607 16450 5616
rect 16500 5630 16620 5658
rect 16408 5370 16436 5607
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 16212 4820 16264 4826
rect 16212 4762 16264 4768
rect 16396 4752 16448 4758
rect 16396 4694 16448 4700
rect 15752 4616 15804 4622
rect 15752 4558 15804 4564
rect 15568 4480 15620 4486
rect 15620 4428 15976 4434
rect 15568 4422 15976 4428
rect 15580 4406 15976 4422
rect 15948 4162 15976 4406
rect 15844 4140 15896 4146
rect 15948 4134 16252 4162
rect 15844 4082 15896 4088
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 15384 2848 15436 2854
rect 15384 2790 15436 2796
rect 15010 2204 15318 2213
rect 15010 2202 15016 2204
rect 15072 2202 15096 2204
rect 15152 2202 15176 2204
rect 15232 2202 15256 2204
rect 15312 2202 15318 2204
rect 15072 2150 15074 2202
rect 15254 2150 15256 2202
rect 15010 2148 15016 2150
rect 15072 2148 15096 2150
rect 15152 2148 15176 2150
rect 15232 2148 15256 2150
rect 15312 2148 15318 2150
rect 15010 2139 15318 2148
rect 14924 740 14976 746
rect 14924 682 14976 688
rect 14832 536 14884 542
rect 14832 478 14884 484
rect 14660 56 14780 82
rect 14844 56 14872 478
rect 15016 264 15068 270
rect 15016 206 15068 212
rect 15028 56 15056 206
rect 15396 56 15424 2790
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 15488 2446 15516 2586
rect 15568 2576 15620 2582
rect 15568 2518 15620 2524
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 15580 56 15608 2518
rect 15672 1562 15700 3878
rect 15752 2848 15804 2854
rect 15752 2790 15804 2796
rect 15660 1556 15712 1562
rect 15660 1498 15712 1504
rect 15764 56 15792 2790
rect 15856 1290 15884 4082
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 15948 2990 15976 3130
rect 16028 3052 16080 3058
rect 16028 2994 16080 3000
rect 15936 2984 15988 2990
rect 15936 2926 15988 2932
rect 16040 2825 16068 2994
rect 16120 2848 16172 2854
rect 16026 2816 16082 2825
rect 16120 2790 16172 2796
rect 16026 2751 16082 2760
rect 15936 2372 15988 2378
rect 15936 2314 15988 2320
rect 15844 1284 15896 1290
rect 15844 1226 15896 1232
rect 15948 56 15976 2314
rect 16132 56 16160 2790
rect 16224 2774 16252 4134
rect 16224 2746 16344 2774
rect 16316 2514 16344 2746
rect 16304 2508 16356 2514
rect 16304 2450 16356 2456
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 16224 2106 16252 2382
rect 16304 2304 16356 2310
rect 16304 2246 16356 2252
rect 16212 2100 16264 2106
rect 16212 2042 16264 2048
rect 16316 56 16344 2246
rect 16408 2106 16436 4694
rect 16500 4486 16528 5630
rect 16960 5234 16988 9279
rect 17144 8634 17172 11096
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17038 8528 17094 8537
rect 17038 8463 17094 8472
rect 17052 5914 17080 8463
rect 17224 8084 17276 8090
rect 17224 8026 17276 8032
rect 17236 7342 17264 8026
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 17328 5098 17356 8910
rect 18708 8634 18736 11096
rect 20272 8634 20300 11096
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17420 8362 17448 8434
rect 17498 8392 17554 8401
rect 17408 8356 17460 8362
rect 17498 8327 17554 8336
rect 19432 8356 19484 8362
rect 17408 8298 17460 8304
rect 17512 5710 17540 8327
rect 19432 8298 19484 8304
rect 18970 7848 19026 7857
rect 17592 7812 17644 7818
rect 18970 7783 19026 7792
rect 19156 7812 19208 7818
rect 17592 7754 17644 7760
rect 17604 7546 17632 7754
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 18052 7404 18104 7410
rect 18052 7346 18104 7352
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17972 5166 18000 7142
rect 18064 6934 18092 7346
rect 18236 7200 18288 7206
rect 18236 7142 18288 7148
rect 18052 6928 18104 6934
rect 18052 6870 18104 6876
rect 18248 5234 18276 7142
rect 18984 6322 19012 7783
rect 19156 7754 19208 7760
rect 19168 6458 19196 7754
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 18984 6118 19012 6258
rect 18972 6112 19024 6118
rect 18972 6054 19024 6060
rect 18236 5228 18288 5234
rect 18236 5170 18288 5176
rect 17960 5160 18012 5166
rect 17960 5102 18012 5108
rect 17316 5092 17368 5098
rect 17316 5034 17368 5040
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 17144 4808 17172 4966
rect 17144 4780 17356 4808
rect 17130 4584 17186 4593
rect 17130 4519 17186 4528
rect 16488 4480 16540 4486
rect 16488 4422 16540 4428
rect 17144 3670 17172 4519
rect 16580 3664 16632 3670
rect 16580 3606 16632 3612
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 16592 2922 16620 3606
rect 16762 3496 16818 3505
rect 16762 3431 16818 3440
rect 16776 3058 16804 3431
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 17224 2984 17276 2990
rect 16960 2932 17224 2938
rect 16960 2926 17276 2932
rect 16580 2916 16632 2922
rect 16580 2858 16632 2864
rect 16960 2910 17264 2926
rect 16672 2848 16724 2854
rect 16672 2790 16724 2796
rect 16488 2576 16540 2582
rect 16488 2518 16540 2524
rect 16396 2100 16448 2106
rect 16396 2042 16448 2048
rect 16500 56 16528 2518
rect 16684 56 16712 2790
rect 16960 2774 16988 2910
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 16776 2746 16988 2774
rect 16776 1737 16804 2746
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 16856 2304 16908 2310
rect 16856 2246 16908 2252
rect 16762 1728 16818 1737
rect 16762 1663 16818 1672
rect 16868 56 16896 2246
rect 16960 1698 16988 2382
rect 16948 1692 17000 1698
rect 16948 1634 17000 1640
rect 17052 56 17080 2790
rect 17328 2774 17356 4780
rect 19248 4548 19300 4554
rect 19248 4490 19300 4496
rect 18972 3732 19024 3738
rect 18972 3674 19024 3680
rect 17776 3528 17828 3534
rect 17828 3488 17908 3516
rect 17776 3470 17828 3476
rect 17408 3460 17460 3466
rect 17408 3402 17460 3408
rect 17500 3460 17552 3466
rect 17500 3402 17552 3408
rect 17420 3058 17448 3402
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 17144 2746 17356 2774
rect 17144 1970 17172 2746
rect 17316 2440 17368 2446
rect 17316 2382 17368 2388
rect 17224 2304 17276 2310
rect 17224 2246 17276 2252
rect 17132 1964 17184 1970
rect 17132 1906 17184 1912
rect 17236 56 17264 2246
rect 17328 1902 17356 2382
rect 17316 1896 17368 1902
rect 17316 1838 17368 1844
rect 17420 56 17448 2790
rect 17512 1873 17540 3402
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 17684 3392 17736 3398
rect 17684 3334 17736 3340
rect 17604 3194 17632 3334
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17592 2304 17644 2310
rect 17592 2246 17644 2252
rect 17498 1864 17554 1873
rect 17498 1799 17554 1808
rect 17604 56 17632 2246
rect 17696 1193 17724 3334
rect 17880 2922 17908 3488
rect 18984 3058 19012 3674
rect 19156 3392 19208 3398
rect 19156 3334 19208 3340
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 17776 2916 17828 2922
rect 17776 2858 17828 2864
rect 17868 2916 17920 2922
rect 17868 2858 17920 2864
rect 19064 2916 19116 2922
rect 19064 2858 19116 2864
rect 17788 2514 17816 2858
rect 18880 2848 18932 2854
rect 18880 2790 18932 2796
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 18144 2576 18196 2582
rect 18144 2518 18196 2524
rect 17776 2508 17828 2514
rect 17776 2450 17828 2456
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 17776 2304 17828 2310
rect 17776 2246 17828 2252
rect 17960 2304 18012 2310
rect 17960 2246 18012 2252
rect 17682 1184 17738 1193
rect 17682 1119 17738 1128
rect 17788 56 17816 2246
rect 17972 56 18000 2246
rect 18064 1766 18092 2382
rect 18052 1760 18104 1766
rect 18052 1702 18104 1708
rect 18156 56 18184 2518
rect 18420 2440 18472 2446
rect 18420 2382 18472 2388
rect 18328 2304 18380 2310
rect 18328 2246 18380 2252
rect 18340 56 18368 2246
rect 18432 2038 18460 2382
rect 18420 2032 18472 2038
rect 18420 1974 18472 1980
rect 18524 56 18552 2586
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 18604 2032 18656 2038
rect 18604 1974 18656 1980
rect 18616 1494 18644 1974
rect 18604 1488 18656 1494
rect 18604 1430 18656 1436
rect 18708 56 18736 2246
rect 18892 56 18920 2790
rect 19076 2514 19104 2858
rect 19064 2508 19116 2514
rect 19064 2450 19116 2456
rect 19064 2372 19116 2378
rect 19064 2314 19116 2320
rect 19076 56 19104 2314
rect 19168 1902 19196 3334
rect 19260 3058 19288 4490
rect 19248 3052 19300 3058
rect 19248 2994 19300 3000
rect 19352 2922 19380 7686
rect 19444 6390 19472 8298
rect 19720 6458 19748 8570
rect 20640 8498 20668 8774
rect 21010 8732 21318 8741
rect 21010 8730 21016 8732
rect 21072 8730 21096 8732
rect 21152 8730 21176 8732
rect 21232 8730 21256 8732
rect 21312 8730 21318 8732
rect 21072 8678 21074 8730
rect 21254 8678 21256 8730
rect 21010 8676 21016 8678
rect 21072 8676 21096 8678
rect 21152 8676 21176 8678
rect 21232 8676 21256 8678
rect 21312 8676 21318 8678
rect 21010 8667 21318 8676
rect 21836 8634 21864 11096
rect 23400 8634 23428 11096
rect 24964 8634 24992 11096
rect 25780 9104 25832 9110
rect 25780 9046 25832 9052
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 23388 8628 23440 8634
rect 23388 8570 23440 8576
rect 24952 8628 25004 8634
rect 24952 8570 25004 8576
rect 25320 8560 25372 8566
rect 25320 8502 25372 8508
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 24860 8492 24912 8498
rect 24860 8434 24912 8440
rect 24768 8288 24820 8294
rect 24768 8230 24820 8236
rect 19950 8188 20258 8197
rect 19950 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20196 8188
rect 20252 8186 20258 8188
rect 20012 8134 20014 8186
rect 20194 8134 20196 8186
rect 19950 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20196 8134
rect 20252 8132 20258 8134
rect 19950 8123 20258 8132
rect 24216 7948 24268 7954
rect 24216 7890 24268 7896
rect 24584 7948 24636 7954
rect 24584 7890 24636 7896
rect 23020 7880 23072 7886
rect 23020 7822 23072 7828
rect 21010 7644 21318 7653
rect 21010 7642 21016 7644
rect 21072 7642 21096 7644
rect 21152 7642 21176 7644
rect 21232 7642 21256 7644
rect 21312 7642 21318 7644
rect 21072 7590 21074 7642
rect 21254 7590 21256 7642
rect 21010 7588 21016 7590
rect 21072 7588 21096 7590
rect 21152 7588 21176 7590
rect 21232 7588 21256 7590
rect 21312 7588 21318 7590
rect 21010 7579 21318 7588
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 21824 7404 21876 7410
rect 21824 7346 21876 7352
rect 19812 6662 19840 7346
rect 19950 7100 20258 7109
rect 19950 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20196 7100
rect 20252 7098 20258 7100
rect 20012 7046 20014 7098
rect 20194 7046 20196 7098
rect 19950 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20196 7046
rect 20252 7044 20258 7046
rect 19950 7035 20258 7044
rect 21836 7002 21864 7346
rect 22008 7200 22060 7206
rect 22008 7142 22060 7148
rect 22284 7200 22336 7206
rect 22284 7142 22336 7148
rect 21824 6996 21876 7002
rect 21824 6938 21876 6944
rect 19800 6656 19852 6662
rect 19800 6598 19852 6604
rect 20444 6656 20496 6662
rect 20444 6598 20496 6604
rect 19708 6452 19760 6458
rect 19708 6394 19760 6400
rect 19432 6384 19484 6390
rect 19432 6326 19484 6332
rect 19950 6012 20258 6021
rect 19950 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20196 6012
rect 20252 6010 20258 6012
rect 20012 5958 20014 6010
rect 20194 5958 20196 6010
rect 19950 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20196 5958
rect 20252 5956 20258 5958
rect 19950 5947 20258 5956
rect 20456 5914 20484 6598
rect 21010 6556 21318 6565
rect 21010 6554 21016 6556
rect 21072 6554 21096 6556
rect 21152 6554 21176 6556
rect 21232 6554 21256 6556
rect 21312 6554 21318 6556
rect 21072 6502 21074 6554
rect 21254 6502 21256 6554
rect 21010 6500 21016 6502
rect 21072 6500 21096 6502
rect 21152 6500 21176 6502
rect 21232 6500 21256 6502
rect 21312 6500 21318 6502
rect 21010 6491 21318 6500
rect 20444 5908 20496 5914
rect 20444 5850 20496 5856
rect 21010 5468 21318 5477
rect 21010 5466 21016 5468
rect 21072 5466 21096 5468
rect 21152 5466 21176 5468
rect 21232 5466 21256 5468
rect 21312 5466 21318 5468
rect 21072 5414 21074 5466
rect 21254 5414 21256 5466
rect 21010 5412 21016 5414
rect 21072 5412 21096 5414
rect 21152 5412 21176 5414
rect 21232 5412 21256 5414
rect 21312 5412 21318 5414
rect 21010 5403 21318 5412
rect 19432 5296 19484 5302
rect 19432 5238 19484 5244
rect 19340 2916 19392 2922
rect 19340 2858 19392 2864
rect 19248 2848 19300 2854
rect 19248 2790 19300 2796
rect 19156 1896 19208 1902
rect 19156 1838 19208 1844
rect 19260 56 19288 2790
rect 19444 2514 19472 5238
rect 21732 5092 21784 5098
rect 21732 5034 21784 5040
rect 19950 4924 20258 4933
rect 19950 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20196 4924
rect 20252 4922 20258 4924
rect 20012 4870 20014 4922
rect 20194 4870 20196 4922
rect 19950 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20196 4870
rect 20252 4868 20258 4870
rect 19950 4859 20258 4868
rect 20810 4720 20866 4729
rect 20628 4684 20680 4690
rect 20810 4655 20866 4664
rect 20628 4626 20680 4632
rect 20444 4276 20496 4282
rect 20444 4218 20496 4224
rect 19950 3836 20258 3845
rect 19950 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20196 3836
rect 20252 3834 20258 3836
rect 20012 3782 20014 3834
rect 20194 3782 20196 3834
rect 19950 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20196 3782
rect 20252 3780 20258 3782
rect 19950 3771 20258 3780
rect 19708 3596 19760 3602
rect 19708 3538 19760 3544
rect 19616 3392 19668 3398
rect 19536 3352 19616 3380
rect 19432 2508 19484 2514
rect 19432 2450 19484 2456
rect 19340 2440 19392 2446
rect 19536 2394 19564 3352
rect 19616 3334 19668 3340
rect 19720 3058 19748 3538
rect 20352 3460 20404 3466
rect 20352 3402 20404 3408
rect 19708 3052 19760 3058
rect 19708 2994 19760 3000
rect 20364 2990 20392 3402
rect 20456 3058 20484 4218
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 20640 2990 20668 4626
rect 20718 3632 20774 3641
rect 20718 3567 20720 3576
rect 20772 3567 20774 3576
rect 20720 3538 20772 3544
rect 20352 2984 20404 2990
rect 20352 2926 20404 2932
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 19708 2916 19760 2922
rect 19708 2858 19760 2864
rect 19800 2916 19852 2922
rect 19800 2858 19852 2864
rect 20536 2916 20588 2922
rect 20536 2858 20588 2864
rect 19616 2848 19668 2854
rect 19616 2790 19668 2796
rect 19340 2382 19392 2388
rect 19352 1834 19380 2382
rect 19444 2366 19564 2394
rect 19340 1828 19392 1834
rect 19340 1770 19392 1776
rect 19444 1465 19472 2366
rect 19524 1488 19576 1494
rect 19430 1456 19486 1465
rect 19524 1430 19576 1436
rect 19430 1391 19486 1400
rect 19536 82 19564 1430
rect 19444 56 19564 82
rect 19628 56 19656 2790
rect 19720 1873 19748 2858
rect 19706 1864 19762 1873
rect 19706 1799 19762 1808
rect 19708 1420 19760 1426
rect 19708 1362 19760 1368
rect 19720 82 19748 1362
rect 19812 218 19840 2858
rect 20352 2848 20404 2854
rect 20352 2790 20404 2796
rect 19950 2748 20258 2757
rect 19950 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20196 2748
rect 20252 2746 20258 2748
rect 20012 2694 20014 2746
rect 20194 2694 20196 2746
rect 19950 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20196 2694
rect 20252 2692 20258 2694
rect 19950 2683 20258 2692
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 19892 2576 19944 2582
rect 19892 2518 19944 2524
rect 19904 1494 19932 2518
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 19996 2106 20024 2382
rect 19984 2100 20036 2106
rect 19984 2042 20036 2048
rect 19892 1488 19944 1494
rect 19892 1430 19944 1436
rect 19812 190 19932 218
rect 19904 82 19932 190
rect 19720 56 19840 82
rect 19904 56 20024 82
rect 20180 56 20208 2586
rect 20260 2304 20312 2310
rect 20260 2246 20312 2252
rect 20272 1426 20300 2246
rect 20260 1420 20312 1426
rect 20260 1362 20312 1368
rect 20364 56 20392 2790
rect 20444 2372 20496 2378
rect 20444 2314 20496 2320
rect 20456 1970 20484 2314
rect 20444 1964 20496 1970
rect 20444 1906 20496 1912
rect 20548 56 20576 2858
rect 20720 2848 20772 2854
rect 20720 2790 20772 2796
rect 20732 56 20760 2790
rect 20824 2446 20852 4655
rect 21010 4380 21318 4389
rect 21010 4378 21016 4380
rect 21072 4378 21096 4380
rect 21152 4378 21176 4380
rect 21232 4378 21256 4380
rect 21312 4378 21318 4380
rect 21072 4326 21074 4378
rect 21254 4326 21256 4378
rect 21010 4324 21016 4326
rect 21072 4324 21096 4326
rect 21152 4324 21176 4326
rect 21232 4324 21256 4326
rect 21312 4324 21318 4326
rect 21010 4315 21318 4324
rect 21364 4208 21416 4214
rect 21364 4150 21416 4156
rect 20904 3664 20956 3670
rect 20904 3606 20956 3612
rect 20916 2774 20944 3606
rect 21010 3292 21318 3301
rect 21010 3290 21016 3292
rect 21072 3290 21096 3292
rect 21152 3290 21176 3292
rect 21232 3290 21256 3292
rect 21312 3290 21318 3292
rect 21072 3238 21074 3290
rect 21254 3238 21256 3290
rect 21010 3236 21016 3238
rect 21072 3236 21096 3238
rect 21152 3236 21176 3238
rect 21232 3236 21256 3238
rect 21312 3236 21318 3238
rect 21010 3227 21318 3236
rect 21376 2938 21404 4150
rect 21640 3392 21692 3398
rect 21638 3360 21640 3369
rect 21692 3360 21694 3369
rect 21638 3295 21694 3304
rect 21284 2910 21404 2938
rect 21640 2916 21692 2922
rect 20916 2746 21036 2774
rect 20904 2576 20956 2582
rect 20904 2518 20956 2524
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 20916 56 20944 2518
rect 21008 2310 21036 2746
rect 21284 2514 21312 2910
rect 21640 2858 21692 2864
rect 21456 2848 21508 2854
rect 21376 2808 21456 2836
rect 21272 2508 21324 2514
rect 21272 2450 21324 2456
rect 20996 2304 21048 2310
rect 20996 2246 21048 2252
rect 21010 2204 21318 2213
rect 21010 2202 21016 2204
rect 21072 2202 21096 2204
rect 21152 2202 21176 2204
rect 21232 2202 21256 2204
rect 21312 2202 21318 2204
rect 21072 2150 21074 2202
rect 21254 2150 21256 2202
rect 21010 2148 21016 2150
rect 21072 2148 21096 2150
rect 21152 2148 21176 2150
rect 21232 2148 21256 2150
rect 21312 2148 21318 2150
rect 21010 2139 21318 2148
rect 21088 1420 21140 1426
rect 21088 1362 21140 1368
rect 21100 56 21128 1362
rect 21376 82 21404 2808
rect 21456 2790 21508 2796
rect 21456 2372 21508 2378
rect 21456 2314 21508 2320
rect 21284 56 21404 82
rect 21468 56 21496 2314
rect 21548 2304 21600 2310
rect 21548 2246 21600 2252
rect 21560 1494 21588 2246
rect 21548 1488 21600 1494
rect 21548 1430 21600 1436
rect 21652 56 21680 2858
rect 21744 2446 21772 5034
rect 22020 4826 22048 7142
rect 22296 5817 22324 7142
rect 22282 5808 22338 5817
rect 22282 5743 22338 5752
rect 22008 4820 22060 4826
rect 22008 4762 22060 4768
rect 22836 4140 22888 4146
rect 22836 4082 22888 4088
rect 21824 4072 21876 4078
rect 21824 4014 21876 4020
rect 21836 3058 21864 4014
rect 22284 4004 22336 4010
rect 22284 3946 22336 3952
rect 21916 3528 21968 3534
rect 21916 3470 21968 3476
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 21824 2644 21876 2650
rect 21824 2586 21876 2592
rect 21732 2440 21784 2446
rect 21732 2382 21784 2388
rect 21732 2304 21784 2310
rect 21732 2246 21784 2252
rect 21744 1426 21772 2246
rect 21732 1420 21784 1426
rect 21732 1362 21784 1368
rect 21836 56 21864 2586
rect 21928 2009 21956 3470
rect 22100 3392 22152 3398
rect 22192 3392 22244 3398
rect 22100 3334 22152 3340
rect 22190 3360 22192 3369
rect 22244 3360 22246 3369
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 21914 2000 21970 2009
rect 21914 1935 21970 1944
rect 22020 56 22048 3130
rect 22112 1970 22140 3334
rect 22190 3295 22246 3304
rect 22296 3058 22324 3946
rect 22376 3596 22428 3602
rect 22376 3538 22428 3544
rect 22284 3052 22336 3058
rect 22284 2994 22336 3000
rect 22192 2576 22244 2582
rect 22192 2518 22244 2524
rect 22100 1964 22152 1970
rect 22100 1906 22152 1912
rect 22204 56 22232 2518
rect 22388 2106 22416 3538
rect 22848 3058 22876 4082
rect 22836 3052 22888 3058
rect 22836 2994 22888 3000
rect 22928 2984 22980 2990
rect 22928 2926 22980 2932
rect 22468 2916 22520 2922
rect 22468 2858 22520 2864
rect 22376 2100 22428 2106
rect 22376 2042 22428 2048
rect 22480 82 22508 2858
rect 22744 2848 22796 2854
rect 22744 2790 22796 2796
rect 22652 2644 22704 2650
rect 22652 2586 22704 2592
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 22572 2038 22600 2382
rect 22560 2032 22612 2038
rect 22560 1974 22612 1980
rect 22664 82 22692 2586
rect 22388 56 22508 82
rect 22572 56 22692 82
rect 22756 56 22784 2790
rect 22940 56 22968 2926
rect 23032 2689 23060 7822
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 24136 6934 24164 7482
rect 24228 7410 24256 7890
rect 24216 7404 24268 7410
rect 24216 7346 24268 7352
rect 24124 6928 24176 6934
rect 24124 6870 24176 6876
rect 24492 6724 24544 6730
rect 24492 6666 24544 6672
rect 24400 6656 24452 6662
rect 24400 6598 24452 6604
rect 24412 6458 24440 6598
rect 24504 6458 24532 6666
rect 24400 6452 24452 6458
rect 24400 6394 24452 6400
rect 24492 6452 24544 6458
rect 24492 6394 24544 6400
rect 24596 6322 24624 7890
rect 24780 7546 24808 8230
rect 24768 7540 24820 7546
rect 24768 7482 24820 7488
rect 24768 7336 24820 7342
rect 24768 7278 24820 7284
rect 24780 7002 24808 7278
rect 24768 6996 24820 7002
rect 24768 6938 24820 6944
rect 24676 6792 24728 6798
rect 24676 6734 24728 6740
rect 24584 6316 24636 6322
rect 24584 6258 24636 6264
rect 23204 4752 23256 4758
rect 23204 4694 23256 4700
rect 23216 3058 23244 4694
rect 24688 4570 24716 6734
rect 24872 6662 24900 8434
rect 24952 8084 25004 8090
rect 24952 8026 25004 8032
rect 24860 6656 24912 6662
rect 24860 6598 24912 6604
rect 24860 5840 24912 5846
rect 24858 5808 24860 5817
rect 24912 5808 24914 5817
rect 24858 5743 24914 5752
rect 24320 4542 24716 4570
rect 23940 4072 23992 4078
rect 23940 4014 23992 4020
rect 23388 3596 23440 3602
rect 23388 3538 23440 3544
rect 23204 3052 23256 3058
rect 23204 2994 23256 3000
rect 23296 2916 23348 2922
rect 23296 2858 23348 2864
rect 23018 2680 23074 2689
rect 23018 2615 23074 2624
rect 23020 2440 23072 2446
rect 23020 2382 23072 2388
rect 23032 1562 23060 2382
rect 23204 2304 23256 2310
rect 23204 2246 23256 2252
rect 23020 1556 23072 1562
rect 23020 1498 23072 1504
rect 23216 82 23244 2246
rect 23124 56 23244 82
rect 23308 56 23336 2858
rect 23400 2553 23428 3538
rect 23572 3392 23624 3398
rect 23572 3334 23624 3340
rect 23584 3097 23612 3334
rect 23664 3188 23716 3194
rect 23664 3130 23716 3136
rect 23570 3088 23626 3097
rect 23570 3023 23626 3032
rect 23480 2576 23532 2582
rect 23386 2544 23442 2553
rect 23480 2518 23532 2524
rect 23386 2479 23442 2488
rect 23492 56 23520 2518
rect 23572 2440 23624 2446
rect 23572 2382 23624 2388
rect 23584 2106 23612 2382
rect 23572 2100 23624 2106
rect 23572 2042 23624 2048
rect 23676 56 23704 3130
rect 23952 3058 23980 4014
rect 24124 3732 24176 3738
rect 24124 3674 24176 3680
rect 24136 3505 24164 3674
rect 24122 3496 24178 3505
rect 24122 3431 24178 3440
rect 23940 3052 23992 3058
rect 23940 2994 23992 3000
rect 24032 2916 24084 2922
rect 24032 2858 24084 2864
rect 23938 2544 23994 2553
rect 23938 2479 23994 2488
rect 23952 2446 23980 2479
rect 23940 2440 23992 2446
rect 23940 2382 23992 2388
rect 23848 2372 23900 2378
rect 23848 2314 23900 2320
rect 23860 56 23888 2314
rect 24044 56 24072 2858
rect 24216 2644 24268 2650
rect 24216 2586 24268 2592
rect 24228 56 24256 2586
rect 24320 1834 24348 4542
rect 24492 4480 24544 4486
rect 24492 4422 24544 4428
rect 24400 2848 24452 2854
rect 24400 2790 24452 2796
rect 24308 1828 24360 1834
rect 24308 1770 24360 1776
rect 24412 56 24440 2790
rect 24504 2446 24532 4422
rect 24676 4004 24728 4010
rect 24676 3946 24728 3952
rect 24584 3392 24636 3398
rect 24584 3334 24636 3340
rect 24596 3097 24624 3334
rect 24582 3088 24638 3097
rect 24688 3058 24716 3946
rect 24768 3664 24820 3670
rect 24766 3632 24768 3641
rect 24820 3632 24822 3641
rect 24766 3567 24822 3576
rect 24860 3528 24912 3534
rect 24860 3470 24912 3476
rect 24768 3188 24820 3194
rect 24768 3130 24820 3136
rect 24582 3023 24638 3032
rect 24676 3052 24728 3058
rect 24676 2994 24728 3000
rect 24492 2440 24544 2446
rect 24492 2382 24544 2388
rect 24584 2304 24636 2310
rect 24584 2246 24636 2252
rect 24596 56 24624 2246
rect 24780 56 24808 3130
rect 24872 2961 24900 3470
rect 24858 2952 24914 2961
rect 24858 2887 24914 2896
rect 24964 2530 24992 8026
rect 25332 7546 25360 8502
rect 25320 7540 25372 7546
rect 25320 7482 25372 7488
rect 25596 7404 25648 7410
rect 25596 7346 25648 7352
rect 25412 6792 25464 6798
rect 25412 6734 25464 6740
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 25148 6390 25176 6598
rect 25136 6384 25188 6390
rect 25136 6326 25188 6332
rect 25136 4616 25188 4622
rect 25136 4558 25188 4564
rect 25044 3460 25096 3466
rect 25044 3402 25096 3408
rect 25056 3058 25084 3402
rect 25044 3052 25096 3058
rect 25044 2994 25096 3000
rect 25148 2904 25176 4558
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 25332 3398 25360 3538
rect 25320 3392 25372 3398
rect 25320 3334 25372 3340
rect 25148 2876 25360 2904
rect 24964 2502 25084 2530
rect 25056 82 25084 2502
rect 25332 2446 25360 2876
rect 25320 2440 25372 2446
rect 25320 2382 25372 2388
rect 25318 1864 25374 1873
rect 25318 1799 25374 1808
rect 24964 56 25084 82
rect 7654 0 7710 40
rect 7838 0 7894 56
rect 8022 0 8078 56
rect 8206 0 8262 56
rect 8390 0 8446 56
rect 8574 0 8630 56
rect 8758 0 8814 56
rect 8864 54 8998 56
rect 8942 0 8998 54
rect 9126 0 9182 56
rect 9310 0 9366 56
rect 9494 0 9550 56
rect 9678 0 9734 56
rect 9862 0 9918 56
rect 10046 0 10102 56
rect 10230 0 10286 56
rect 10414 0 10470 56
rect 10598 0 10654 56
rect 10782 0 10838 56
rect 10966 0 11022 56
rect 11150 0 11206 56
rect 11334 0 11390 56
rect 11518 0 11574 56
rect 11702 0 11758 56
rect 11886 54 12020 56
rect 11886 0 11942 54
rect 12070 0 12126 56
rect 12254 0 12310 56
rect 12438 0 12494 56
rect 12622 0 12678 56
rect 12806 0 12862 56
rect 12990 0 13046 56
rect 13174 0 13230 56
rect 13358 0 13414 56
rect 13542 0 13598 56
rect 13726 0 13782 56
rect 13910 0 13966 56
rect 14094 54 14228 56
rect 14278 54 14412 56
rect 14094 0 14150 54
rect 14278 0 14334 54
rect 14462 0 14518 56
rect 14646 54 14780 56
rect 14646 0 14702 54
rect 14830 0 14886 56
rect 15014 0 15070 56
rect 15198 0 15254 56
rect 15382 0 15438 56
rect 15566 0 15622 56
rect 15750 0 15806 56
rect 15934 0 15990 56
rect 16118 0 16174 56
rect 16302 0 16358 56
rect 16486 0 16542 56
rect 16670 0 16726 56
rect 16854 0 16910 56
rect 17038 0 17094 56
rect 17222 0 17278 56
rect 17406 0 17462 56
rect 17590 0 17646 56
rect 17774 0 17830 56
rect 17958 0 18014 56
rect 18142 0 18198 56
rect 18326 0 18382 56
rect 18510 0 18566 56
rect 18694 0 18750 56
rect 18878 0 18934 56
rect 19062 0 19118 56
rect 19246 0 19302 56
rect 19430 54 19564 56
rect 19430 0 19486 54
rect 19614 0 19670 56
rect 19720 54 19854 56
rect 19904 54 20038 56
rect 19798 0 19854 54
rect 19982 0 20038 54
rect 20166 0 20222 56
rect 20350 0 20406 56
rect 20534 0 20590 56
rect 20718 0 20774 56
rect 20902 0 20958 56
rect 21086 0 21142 56
rect 21270 54 21404 56
rect 21270 0 21326 54
rect 21454 0 21510 56
rect 21638 0 21694 56
rect 21822 0 21878 56
rect 22006 0 22062 56
rect 22190 0 22246 56
rect 22374 54 22508 56
rect 22558 54 22692 56
rect 22374 0 22430 54
rect 22558 0 22614 54
rect 22742 0 22798 56
rect 22926 0 22982 56
rect 23110 54 23244 56
rect 23110 0 23166 54
rect 23294 0 23350 56
rect 23478 0 23534 56
rect 23662 0 23718 56
rect 23846 0 23902 56
rect 24030 0 24086 56
rect 24214 0 24270 56
rect 24398 0 24454 56
rect 24582 0 24638 56
rect 24766 0 24822 56
rect 24950 54 25084 56
rect 25134 96 25190 105
rect 24950 0 25006 54
rect 25332 56 25360 1799
rect 25424 105 25452 6734
rect 25504 3936 25556 3942
rect 25504 3878 25556 3884
rect 25516 3058 25544 3878
rect 25504 3052 25556 3058
rect 25504 2994 25556 3000
rect 25502 2680 25558 2689
rect 25502 2615 25558 2624
rect 25516 898 25544 2615
rect 25608 1329 25636 7346
rect 25688 7336 25740 7342
rect 25688 7278 25740 7284
rect 25594 1320 25650 1329
rect 25594 1255 25650 1264
rect 25516 870 25636 898
rect 25504 740 25556 746
rect 25504 682 25556 688
rect 25410 96 25466 105
rect 25134 0 25190 40
rect 25318 0 25374 56
rect 25516 56 25544 682
rect 25608 82 25636 870
rect 25700 762 25728 7278
rect 25792 6662 25820 9046
rect 26528 8634 26556 11096
rect 27436 8832 27488 8838
rect 27436 8774 27488 8780
rect 27010 8732 27318 8741
rect 27010 8730 27016 8732
rect 27072 8730 27096 8732
rect 27152 8730 27176 8732
rect 27232 8730 27256 8732
rect 27312 8730 27318 8732
rect 27072 8678 27074 8730
rect 27254 8678 27256 8730
rect 27010 8676 27016 8678
rect 27072 8676 27096 8678
rect 27152 8676 27176 8678
rect 27232 8676 27256 8678
rect 27312 8676 27318 8678
rect 27010 8667 27318 8676
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 25950 8188 26258 8197
rect 25950 8186 25956 8188
rect 26012 8186 26036 8188
rect 26092 8186 26116 8188
rect 26172 8186 26196 8188
rect 26252 8186 26258 8188
rect 26012 8134 26014 8186
rect 26194 8134 26196 8186
rect 25950 8132 25956 8134
rect 26012 8132 26036 8134
rect 26092 8132 26116 8134
rect 26172 8132 26196 8134
rect 26252 8132 26258 8134
rect 25950 8123 26258 8132
rect 27010 7644 27318 7653
rect 27010 7642 27016 7644
rect 27072 7642 27096 7644
rect 27152 7642 27176 7644
rect 27232 7642 27256 7644
rect 27312 7642 27318 7644
rect 27072 7590 27074 7642
rect 27254 7590 27256 7642
rect 27010 7588 27016 7590
rect 27072 7588 27096 7590
rect 27152 7588 27176 7590
rect 27232 7588 27256 7590
rect 27312 7588 27318 7590
rect 27010 7579 27318 7588
rect 27448 7546 27476 8774
rect 28092 8634 28120 11096
rect 28540 9036 28592 9042
rect 28540 8978 28592 8984
rect 28264 8900 28316 8906
rect 28264 8842 28316 8848
rect 28080 8628 28132 8634
rect 28080 8570 28132 8576
rect 27988 8492 28040 8498
rect 27988 8434 28040 8440
rect 28000 7546 28028 8434
rect 28276 7546 28304 8842
rect 28552 7546 28580 8978
rect 29656 8634 29684 11096
rect 31114 9344 31170 9353
rect 31114 9279 31170 9288
rect 30932 8968 30984 8974
rect 30932 8910 30984 8916
rect 29644 8628 29696 8634
rect 29644 8570 29696 8576
rect 30656 8560 30708 8566
rect 30656 8502 30708 8508
rect 28724 8492 28776 8498
rect 28724 8434 28776 8440
rect 29736 8492 29788 8498
rect 29736 8434 29788 8440
rect 27436 7540 27488 7546
rect 27436 7482 27488 7488
rect 27988 7540 28040 7546
rect 27988 7482 28040 7488
rect 28264 7540 28316 7546
rect 28264 7482 28316 7488
rect 28540 7540 28592 7546
rect 28540 7482 28592 7488
rect 26884 7472 26936 7478
rect 26884 7414 26936 7420
rect 26792 7336 26844 7342
rect 26792 7278 26844 7284
rect 25872 7268 25924 7274
rect 25872 7210 25924 7216
rect 25780 6656 25832 6662
rect 25780 6598 25832 6604
rect 25884 5778 25912 7210
rect 25950 7100 26258 7109
rect 25950 7098 25956 7100
rect 26012 7098 26036 7100
rect 26092 7098 26116 7100
rect 26172 7098 26196 7100
rect 26252 7098 26258 7100
rect 26012 7046 26014 7098
rect 26194 7046 26196 7098
rect 25950 7044 25956 7046
rect 26012 7044 26036 7046
rect 26092 7044 26116 7046
rect 26172 7044 26196 7046
rect 26252 7044 26258 7046
rect 25950 7035 26258 7044
rect 26424 6792 26476 6798
rect 26424 6734 26476 6740
rect 25950 6012 26258 6021
rect 25950 6010 25956 6012
rect 26012 6010 26036 6012
rect 26092 6010 26116 6012
rect 26172 6010 26196 6012
rect 26252 6010 26258 6012
rect 26012 5958 26014 6010
rect 26194 5958 26196 6010
rect 25950 5956 25956 5958
rect 26012 5956 26036 5958
rect 26092 5956 26116 5958
rect 26172 5956 26196 5958
rect 26252 5956 26258 5958
rect 25950 5947 26258 5956
rect 25872 5772 25924 5778
rect 25872 5714 25924 5720
rect 25950 4924 26258 4933
rect 25950 4922 25956 4924
rect 26012 4922 26036 4924
rect 26092 4922 26116 4924
rect 26172 4922 26196 4924
rect 26252 4922 26258 4924
rect 26012 4870 26014 4922
rect 26194 4870 26196 4922
rect 25950 4868 25956 4870
rect 26012 4868 26036 4870
rect 26092 4868 26116 4870
rect 26172 4868 26196 4870
rect 26252 4868 26258 4870
rect 25950 4859 26258 4868
rect 25950 3836 26258 3845
rect 25950 3834 25956 3836
rect 26012 3834 26036 3836
rect 26092 3834 26116 3836
rect 26172 3834 26196 3836
rect 26252 3834 26258 3836
rect 26012 3782 26014 3834
rect 26194 3782 26196 3834
rect 25950 3780 25956 3782
rect 26012 3780 26036 3782
rect 26092 3780 26116 3782
rect 26172 3780 26196 3782
rect 26252 3780 26258 3782
rect 25950 3771 26258 3780
rect 26330 3768 26386 3777
rect 26056 3732 26108 3738
rect 26330 3703 26386 3712
rect 26056 3674 26108 3680
rect 25780 3392 25832 3398
rect 25780 3334 25832 3340
rect 25792 3058 25820 3334
rect 26068 3074 26096 3674
rect 26344 3618 26372 3703
rect 26160 3602 26372 3618
rect 26148 3596 26372 3602
rect 26200 3590 26372 3596
rect 26148 3538 26200 3544
rect 26332 3528 26384 3534
rect 26332 3470 26384 3476
rect 25780 3052 25832 3058
rect 25780 2994 25832 3000
rect 25884 3046 26096 3074
rect 25780 2848 25832 2854
rect 25780 2790 25832 2796
rect 25792 2553 25820 2790
rect 25884 2650 25912 3046
rect 25950 2748 26258 2757
rect 25950 2746 25956 2748
rect 26012 2746 26036 2748
rect 26092 2746 26116 2748
rect 26172 2746 26196 2748
rect 26252 2746 26258 2748
rect 26012 2694 26014 2746
rect 26194 2694 26196 2746
rect 25950 2692 25956 2694
rect 26012 2692 26036 2694
rect 26092 2692 26116 2694
rect 26172 2692 26196 2694
rect 26252 2692 26258 2694
rect 25950 2683 26258 2692
rect 25872 2644 25924 2650
rect 25872 2586 25924 2592
rect 25778 2544 25834 2553
rect 25778 2479 25834 2488
rect 26054 2544 26110 2553
rect 26054 2479 26110 2488
rect 25700 734 25912 762
rect 25608 56 25728 82
rect 25884 56 25912 734
rect 26068 56 26096 2479
rect 26344 82 26372 3470
rect 26252 56 26372 82
rect 26436 56 26464 6734
rect 26608 6724 26660 6730
rect 26608 6666 26660 6672
rect 26700 6724 26752 6730
rect 26700 6666 26752 6672
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 26528 406 26556 3470
rect 26620 1408 26648 6666
rect 26712 5273 26740 6666
rect 26698 5264 26754 5273
rect 26698 5199 26754 5208
rect 26804 3602 26832 7278
rect 26896 3738 26924 7414
rect 27620 7404 27672 7410
rect 27620 7346 27672 7352
rect 27988 7404 28040 7410
rect 27988 7346 28040 7352
rect 28448 7404 28500 7410
rect 28448 7346 28500 7352
rect 27010 6556 27318 6565
rect 27010 6554 27016 6556
rect 27072 6554 27096 6556
rect 27152 6554 27176 6556
rect 27232 6554 27256 6556
rect 27312 6554 27318 6556
rect 27072 6502 27074 6554
rect 27254 6502 27256 6554
rect 27010 6500 27016 6502
rect 27072 6500 27096 6502
rect 27152 6500 27176 6502
rect 27232 6500 27256 6502
rect 27312 6500 27318 6502
rect 27010 6491 27318 6500
rect 27010 5468 27318 5477
rect 27010 5466 27016 5468
rect 27072 5466 27096 5468
rect 27152 5466 27176 5468
rect 27232 5466 27256 5468
rect 27312 5466 27318 5468
rect 27072 5414 27074 5466
rect 27254 5414 27256 5466
rect 27010 5412 27016 5414
rect 27072 5412 27096 5414
rect 27152 5412 27176 5414
rect 27232 5412 27256 5414
rect 27312 5412 27318 5414
rect 27010 5403 27318 5412
rect 27528 4548 27580 4554
rect 27528 4490 27580 4496
rect 27010 4380 27318 4389
rect 27010 4378 27016 4380
rect 27072 4378 27096 4380
rect 27152 4378 27176 4380
rect 27232 4378 27256 4380
rect 27312 4378 27318 4380
rect 27072 4326 27074 4378
rect 27254 4326 27256 4378
rect 27010 4324 27016 4326
rect 27072 4324 27096 4326
rect 27152 4324 27176 4326
rect 27232 4324 27256 4326
rect 27312 4324 27318 4326
rect 27010 4315 27318 4324
rect 27540 4185 27568 4490
rect 27526 4176 27582 4185
rect 27344 4140 27396 4146
rect 27526 4111 27582 4120
rect 27344 4082 27396 4088
rect 26884 3732 26936 3738
rect 26884 3674 26936 3680
rect 26792 3596 26844 3602
rect 26792 3538 26844 3544
rect 26884 3528 26936 3534
rect 26884 3470 26936 3476
rect 26700 3392 26752 3398
rect 26700 3334 26752 3340
rect 26792 3392 26844 3398
rect 26792 3334 26844 3340
rect 26712 2446 26740 3334
rect 26804 2514 26832 3334
rect 26792 2508 26844 2514
rect 26792 2450 26844 2456
rect 26700 2440 26752 2446
rect 26896 2417 26924 3470
rect 27010 3292 27318 3301
rect 27010 3290 27016 3292
rect 27072 3290 27096 3292
rect 27152 3290 27176 3292
rect 27232 3290 27256 3292
rect 27312 3290 27318 3292
rect 27072 3238 27074 3290
rect 27254 3238 27256 3290
rect 27010 3236 27016 3238
rect 27072 3236 27096 3238
rect 27152 3236 27176 3238
rect 27232 3236 27256 3238
rect 27312 3236 27318 3238
rect 27010 3227 27318 3236
rect 27068 3188 27120 3194
rect 27068 3130 27120 3136
rect 26700 2382 26752 2388
rect 26882 2408 26938 2417
rect 26882 2343 26938 2352
rect 27080 2292 27108 3130
rect 26896 2264 27108 2292
rect 26620 1380 26832 1408
rect 26516 400 26568 406
rect 26516 342 26568 348
rect 26606 96 26662 105
rect 25410 31 25466 40
rect 25502 0 25558 56
rect 25608 54 25742 56
rect 25686 0 25742 54
rect 25870 0 25926 56
rect 26054 0 26110 56
rect 26238 54 26372 56
rect 26238 0 26294 54
rect 26422 0 26478 56
rect 26804 56 26832 1380
rect 26896 377 26924 2264
rect 27010 2204 27318 2213
rect 27010 2202 27016 2204
rect 27072 2202 27096 2204
rect 27152 2202 27176 2204
rect 27232 2202 27256 2204
rect 27312 2202 27318 2204
rect 27072 2150 27074 2202
rect 27254 2150 27256 2202
rect 27010 2148 27016 2150
rect 27072 2148 27096 2150
rect 27152 2148 27176 2150
rect 27232 2148 27256 2150
rect 27312 2148 27318 2150
rect 27010 2139 27318 2148
rect 27356 1714 27384 4082
rect 27528 3936 27580 3942
rect 27528 3878 27580 3884
rect 27436 3528 27488 3534
rect 27436 3470 27488 3476
rect 27264 1686 27384 1714
rect 27160 1420 27212 1426
rect 27160 1362 27212 1368
rect 26974 1320 27030 1329
rect 26974 1255 27030 1264
rect 26882 368 26938 377
rect 26882 303 26938 312
rect 26988 56 27016 1255
rect 27172 56 27200 1362
rect 27264 202 27292 1686
rect 27344 1624 27396 1630
rect 27344 1566 27396 1572
rect 27252 196 27304 202
rect 27252 138 27304 144
rect 27356 56 27384 1566
rect 27448 134 27476 3470
rect 27540 3194 27568 3878
rect 27528 3188 27580 3194
rect 27528 3130 27580 3136
rect 27526 1456 27582 1465
rect 27632 1426 27660 7346
rect 27804 4616 27856 4622
rect 27804 4558 27856 4564
rect 27896 4616 27948 4622
rect 27896 4558 27948 4564
rect 27816 4486 27844 4558
rect 27804 4480 27856 4486
rect 27804 4422 27856 4428
rect 27908 4185 27936 4558
rect 27894 4176 27950 4185
rect 27894 4111 27950 4120
rect 27896 4072 27948 4078
rect 27896 4014 27948 4020
rect 27908 3942 27936 4014
rect 27712 3936 27764 3942
rect 27712 3878 27764 3884
rect 27896 3936 27948 3942
rect 27896 3878 27948 3884
rect 27724 2666 27752 3878
rect 27804 3596 27856 3602
rect 27804 3538 27856 3544
rect 27816 3194 27844 3538
rect 27896 3528 27948 3534
rect 27896 3470 27948 3476
rect 27804 3188 27856 3194
rect 27804 3130 27856 3136
rect 27804 3052 27856 3058
rect 27804 2994 27856 3000
rect 27816 2961 27844 2994
rect 27802 2952 27858 2961
rect 27802 2887 27858 2896
rect 27724 2638 27844 2666
rect 27816 2582 27844 2638
rect 27804 2576 27856 2582
rect 27804 2518 27856 2524
rect 27712 1828 27764 1834
rect 27712 1770 27764 1776
rect 27526 1391 27582 1400
rect 27620 1420 27672 1426
rect 27436 128 27488 134
rect 27436 70 27488 76
rect 27540 56 27568 1391
rect 27620 1362 27672 1368
rect 27724 56 27752 1770
rect 27908 354 27936 3470
rect 27816 326 27936 354
rect 27816 134 27844 326
rect 27804 128 27856 134
rect 28000 82 28028 7346
rect 28080 6792 28132 6798
rect 28080 6734 28132 6740
rect 27804 70 27856 76
rect 27908 56 28028 82
rect 28092 56 28120 6734
rect 28460 4729 28488 7346
rect 28736 6662 28764 8434
rect 29460 8356 29512 8362
rect 29460 8298 29512 8304
rect 29472 7546 29500 8298
rect 29460 7540 29512 7546
rect 29460 7482 29512 7488
rect 29644 7404 29696 7410
rect 29644 7346 29696 7352
rect 28724 6656 28776 6662
rect 28724 6598 28776 6604
rect 28632 5228 28684 5234
rect 28632 5170 28684 5176
rect 28446 4720 28502 4729
rect 28446 4655 28502 4664
rect 28264 4616 28316 4622
rect 28262 4584 28264 4593
rect 28316 4584 28318 4593
rect 28262 4519 28318 4528
rect 28448 4072 28500 4078
rect 28446 4040 28448 4049
rect 28500 4040 28502 4049
rect 28446 3975 28502 3984
rect 28356 3528 28408 3534
rect 28262 3496 28318 3505
rect 28356 3470 28408 3476
rect 28262 3431 28318 3440
rect 28172 3392 28224 3398
rect 28172 3334 28224 3340
rect 28184 2106 28212 3334
rect 28276 2922 28304 3431
rect 28264 2916 28316 2922
rect 28264 2858 28316 2864
rect 28172 2100 28224 2106
rect 28172 2042 28224 2048
rect 28264 1420 28316 1426
rect 28264 1362 28316 1368
rect 28276 56 28304 1362
rect 28368 474 28396 3470
rect 28540 3392 28592 3398
rect 28540 3334 28592 3340
rect 28448 3120 28500 3126
rect 28446 3088 28448 3097
rect 28500 3088 28502 3097
rect 28446 3023 28502 3032
rect 28448 1556 28500 1562
rect 28448 1498 28500 1504
rect 28356 468 28408 474
rect 28356 410 28408 416
rect 28460 56 28488 1498
rect 28552 542 28580 3334
rect 28540 536 28592 542
rect 28540 478 28592 484
rect 28644 56 28672 5170
rect 29552 4140 29604 4146
rect 29552 4082 29604 4088
rect 28908 4072 28960 4078
rect 28908 4014 28960 4020
rect 28724 4004 28776 4010
rect 28724 3946 28776 3952
rect 28736 338 28764 3946
rect 28816 3936 28868 3942
rect 28816 3878 28868 3884
rect 28828 2854 28856 3878
rect 28920 3738 28948 4014
rect 29184 3936 29236 3942
rect 29184 3878 29236 3884
rect 28908 3732 28960 3738
rect 28908 3674 28960 3680
rect 28816 2848 28868 2854
rect 28816 2790 28868 2796
rect 29196 1698 29224 3878
rect 29184 1692 29236 1698
rect 29184 1634 29236 1640
rect 28724 332 28776 338
rect 28724 274 28776 280
rect 29564 270 29592 4082
rect 29656 1630 29684 7346
rect 29748 6458 29776 8434
rect 30472 7404 30524 7410
rect 30472 7346 30524 7352
rect 30380 7336 30432 7342
rect 30380 7278 30432 7284
rect 30392 6866 30420 7278
rect 30380 6860 30432 6866
rect 30380 6802 30432 6808
rect 29736 6452 29788 6458
rect 29736 6394 29788 6400
rect 29920 6316 29972 6322
rect 29920 6258 29972 6264
rect 29644 1624 29696 1630
rect 29644 1566 29696 1572
rect 29932 1426 29960 6258
rect 30378 3632 30434 3641
rect 30378 3567 30380 3576
rect 30432 3567 30434 3576
rect 30380 3538 30432 3544
rect 30484 1465 30512 7346
rect 30564 7200 30616 7206
rect 30564 7142 30616 7148
rect 30576 4146 30604 7142
rect 30668 5914 30696 8502
rect 30944 8498 30972 8910
rect 31128 8634 31156 9279
rect 31220 8634 31248 11096
rect 31390 9616 31446 9625
rect 31390 9551 31446 9560
rect 31116 8628 31168 8634
rect 31116 8570 31168 8576
rect 31208 8628 31260 8634
rect 31208 8570 31260 8576
rect 30932 8492 30984 8498
rect 30932 8434 30984 8440
rect 31300 8492 31352 8498
rect 31300 8434 31352 8440
rect 30840 8424 30892 8430
rect 30840 8366 30892 8372
rect 31024 8424 31076 8430
rect 31024 8366 31076 8372
rect 30852 7546 30880 8366
rect 30840 7540 30892 7546
rect 30840 7482 30892 7488
rect 30932 6928 30984 6934
rect 30932 6870 30984 6876
rect 30656 5908 30708 5914
rect 30656 5850 30708 5856
rect 30944 5710 30972 6870
rect 31036 6254 31064 8366
rect 31208 7880 31260 7886
rect 31208 7822 31260 7828
rect 31220 6390 31248 7822
rect 31208 6384 31260 6390
rect 31208 6326 31260 6332
rect 31024 6248 31076 6254
rect 31024 6190 31076 6196
rect 31312 5914 31340 8434
rect 31404 8090 31432 9551
rect 31758 9072 31814 9081
rect 31758 9007 31814 9016
rect 31772 8090 31800 9007
rect 32784 8634 32812 11096
rect 33414 8800 33470 8809
rect 33010 8732 33318 8741
rect 33414 8735 33470 8744
rect 33010 8730 33016 8732
rect 33072 8730 33096 8732
rect 33152 8730 33176 8732
rect 33232 8730 33256 8732
rect 33312 8730 33318 8732
rect 33072 8678 33074 8730
rect 33254 8678 33256 8730
rect 33010 8676 33016 8678
rect 33072 8676 33096 8678
rect 33152 8676 33176 8678
rect 33232 8676 33256 8678
rect 33312 8676 33318 8678
rect 33010 8667 33318 8676
rect 32772 8628 32824 8634
rect 32772 8570 32824 8576
rect 32310 8528 32366 8537
rect 32310 8463 32366 8472
rect 32404 8492 32456 8498
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 32324 8090 32352 8463
rect 32404 8434 32456 8440
rect 31392 8084 31444 8090
rect 31392 8026 31444 8032
rect 31760 8084 31812 8090
rect 31760 8026 31812 8032
rect 32312 8084 32364 8090
rect 32312 8026 32364 8032
rect 31668 7880 31720 7886
rect 31668 7822 31720 7828
rect 31392 7404 31444 7410
rect 31392 7346 31444 7352
rect 31300 5908 31352 5914
rect 31300 5850 31352 5856
rect 30840 5704 30892 5710
rect 30840 5646 30892 5652
rect 30932 5704 30984 5710
rect 30932 5646 30984 5652
rect 30564 4140 30616 4146
rect 30564 4082 30616 4088
rect 30852 1562 30880 5646
rect 31404 5574 31432 7346
rect 31680 5642 31708 7822
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 31852 6996 31904 7002
rect 31852 6938 31904 6944
rect 31760 6792 31812 6798
rect 31760 6734 31812 6740
rect 31668 5636 31720 5642
rect 31668 5578 31720 5584
rect 31392 5568 31444 5574
rect 31392 5510 31444 5516
rect 31772 4690 31800 6734
rect 31760 4684 31812 4690
rect 31760 4626 31812 4632
rect 31864 4622 31892 6938
rect 32312 6316 32364 6322
rect 32312 6258 32364 6264
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 32324 5370 32352 6258
rect 32312 5364 32364 5370
rect 32312 5306 32364 5312
rect 32416 5098 32444 8434
rect 33048 8356 33100 8362
rect 33048 8298 33100 8304
rect 32496 8288 32548 8294
rect 33060 8265 33088 8298
rect 32496 8230 32548 8236
rect 33046 8256 33102 8265
rect 32508 7993 32536 8230
rect 33046 8191 33102 8200
rect 32494 7984 32550 7993
rect 32494 7919 32550 7928
rect 32496 7744 32548 7750
rect 32496 7686 32548 7692
rect 32508 7449 32536 7686
rect 33010 7644 33318 7653
rect 33010 7642 33016 7644
rect 33072 7642 33096 7644
rect 33152 7642 33176 7644
rect 33232 7642 33256 7644
rect 33312 7642 33318 7644
rect 33072 7590 33074 7642
rect 33254 7590 33256 7642
rect 33010 7588 33016 7590
rect 33072 7588 33096 7590
rect 33152 7588 33176 7590
rect 33232 7588 33256 7590
rect 33312 7588 33318 7590
rect 33010 7579 33318 7588
rect 33428 7546 33456 8735
rect 33600 7744 33652 7750
rect 33598 7712 33600 7721
rect 33652 7712 33654 7721
rect 33598 7647 33654 7656
rect 33416 7540 33468 7546
rect 33416 7482 33468 7488
rect 32494 7440 32550 7449
rect 32494 7375 32550 7384
rect 32864 7200 32916 7206
rect 32862 7168 32864 7177
rect 32916 7168 32918 7177
rect 32862 7103 32918 7112
rect 32862 6896 32918 6905
rect 32862 6831 32918 6840
rect 32876 6662 32904 6831
rect 33416 6724 33468 6730
rect 33416 6666 33468 6672
rect 32864 6656 32916 6662
rect 33428 6633 33456 6666
rect 32864 6598 32916 6604
rect 33414 6624 33470 6633
rect 33010 6556 33318 6565
rect 33414 6559 33470 6568
rect 33010 6554 33016 6556
rect 33072 6554 33096 6556
rect 33152 6554 33176 6556
rect 33232 6554 33256 6556
rect 33312 6554 33318 6556
rect 33072 6502 33074 6554
rect 33254 6502 33256 6554
rect 33010 6500 33016 6502
rect 33072 6500 33096 6502
rect 33152 6500 33176 6502
rect 33232 6500 33256 6502
rect 33312 6500 33318 6502
rect 33010 6491 33318 6500
rect 32864 6452 32916 6458
rect 32864 6394 32916 6400
rect 32876 6361 32904 6394
rect 32862 6352 32918 6361
rect 32862 6287 32918 6296
rect 32496 6112 32548 6118
rect 32494 6080 32496 6089
rect 32548 6080 32550 6089
rect 32494 6015 32550 6024
rect 32864 5840 32916 5846
rect 32862 5808 32864 5817
rect 32916 5808 32918 5817
rect 32862 5743 32918 5752
rect 33416 5568 33468 5574
rect 33414 5536 33416 5545
rect 33468 5536 33470 5545
rect 33010 5468 33318 5477
rect 33414 5471 33470 5480
rect 33010 5466 33016 5468
rect 33072 5466 33096 5468
rect 33152 5466 33176 5468
rect 33232 5466 33256 5468
rect 33312 5466 33318 5468
rect 33072 5414 33074 5466
rect 33254 5414 33256 5466
rect 33010 5412 33016 5414
rect 33072 5412 33096 5414
rect 33152 5412 33176 5414
rect 33232 5412 33256 5414
rect 33312 5412 33318 5414
rect 33010 5403 33318 5412
rect 32864 5364 32916 5370
rect 32864 5306 32916 5312
rect 32876 5273 32904 5306
rect 32862 5264 32918 5273
rect 32862 5199 32918 5208
rect 32404 5092 32456 5098
rect 32404 5034 32456 5040
rect 32496 5024 32548 5030
rect 32494 4992 32496 5001
rect 32548 4992 32550 5001
rect 31950 4924 32258 4933
rect 32494 4927 32550 4936
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 32864 4752 32916 4758
rect 32862 4720 32864 4729
rect 32916 4720 32918 4729
rect 32862 4655 32918 4664
rect 31852 4616 31904 4622
rect 31852 4558 31904 4564
rect 33416 4480 33468 4486
rect 33414 4448 33416 4457
rect 33468 4448 33470 4457
rect 33010 4380 33318 4389
rect 33414 4383 33470 4392
rect 33010 4378 33016 4380
rect 33072 4378 33096 4380
rect 33152 4378 33176 4380
rect 33232 4378 33256 4380
rect 33312 4378 33318 4380
rect 33072 4326 33074 4378
rect 33254 4326 33256 4378
rect 33010 4324 33016 4326
rect 33072 4324 33096 4326
rect 33152 4324 33176 4326
rect 33232 4324 33256 4326
rect 33312 4324 33318 4326
rect 33010 4315 33318 4324
rect 32862 4176 32918 4185
rect 32862 4111 32918 4120
rect 32876 4010 32904 4111
rect 32864 4004 32916 4010
rect 32864 3946 32916 3952
rect 32496 3936 32548 3942
rect 32494 3904 32496 3913
rect 32548 3904 32550 3913
rect 31950 3836 32258 3845
rect 32494 3839 32550 3848
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31666 3768 31722 3777
rect 31950 3771 32258 3780
rect 31666 3703 31722 3712
rect 31680 3058 31708 3703
rect 32864 3664 32916 3670
rect 32862 3632 32864 3641
rect 32916 3632 32918 3641
rect 32862 3567 32918 3576
rect 33416 3392 33468 3398
rect 33414 3360 33416 3369
rect 33468 3360 33470 3369
rect 33010 3292 33318 3301
rect 33414 3295 33470 3304
rect 33010 3290 33016 3292
rect 33072 3290 33096 3292
rect 33152 3290 33176 3292
rect 33232 3290 33256 3292
rect 33312 3290 33318 3292
rect 33072 3238 33074 3290
rect 33254 3238 33256 3290
rect 33010 3236 33016 3238
rect 33072 3236 33096 3238
rect 33152 3236 33176 3238
rect 33232 3236 33256 3238
rect 33312 3236 33318 3238
rect 33010 3227 33318 3236
rect 32864 3188 32916 3194
rect 32864 3130 32916 3136
rect 32876 3097 32904 3130
rect 32862 3088 32918 3097
rect 31668 3052 31720 3058
rect 32862 3023 32918 3032
rect 31668 2994 31720 3000
rect 32404 2848 32456 2854
rect 32496 2848 32548 2854
rect 32404 2790 32456 2796
rect 32494 2816 32496 2825
rect 32548 2816 32550 2825
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 30932 2440 30984 2446
rect 30932 2382 30984 2388
rect 31300 2440 31352 2446
rect 31300 2382 31352 2388
rect 31668 2440 31720 2446
rect 31668 2382 31720 2388
rect 32312 2440 32364 2446
rect 32312 2382 32364 2388
rect 30944 1970 30972 2382
rect 31116 2304 31168 2310
rect 31116 2246 31168 2252
rect 31128 2009 31156 2246
rect 31312 2038 31340 2382
rect 31484 2304 31536 2310
rect 31484 2246 31536 2252
rect 31300 2032 31352 2038
rect 31114 2000 31170 2009
rect 30932 1964 30984 1970
rect 31300 1974 31352 1980
rect 31114 1935 31170 1944
rect 30932 1906 30984 1912
rect 30840 1556 30892 1562
rect 30840 1498 30892 1504
rect 31496 1465 31524 2246
rect 31680 1902 31708 2382
rect 31852 2304 31904 2310
rect 31852 2246 31904 2252
rect 31668 1896 31720 1902
rect 31668 1838 31720 1844
rect 30470 1456 30526 1465
rect 29920 1420 29972 1426
rect 30470 1391 30526 1400
rect 31482 1456 31538 1465
rect 31482 1391 31538 1400
rect 29920 1362 29972 1368
rect 31864 1193 31892 2246
rect 32324 1494 32352 2382
rect 32416 1737 32444 2790
rect 32494 2751 32550 2760
rect 32864 2576 32916 2582
rect 32862 2544 32864 2553
rect 32916 2544 32918 2553
rect 32862 2479 32918 2488
rect 33416 2304 33468 2310
rect 33414 2272 33416 2281
rect 33468 2272 33470 2281
rect 33010 2204 33318 2213
rect 33414 2207 33470 2216
rect 33010 2202 33016 2204
rect 33072 2202 33096 2204
rect 33152 2202 33176 2204
rect 33232 2202 33256 2204
rect 33312 2202 33318 2204
rect 33072 2150 33074 2202
rect 33254 2150 33256 2202
rect 33010 2148 33016 2150
rect 33072 2148 33096 2150
rect 33152 2148 33176 2150
rect 33232 2148 33256 2150
rect 33312 2148 33318 2150
rect 33010 2139 33318 2148
rect 32402 1728 32458 1737
rect 32402 1663 32458 1672
rect 32312 1488 32364 1494
rect 32312 1430 32364 1436
rect 31850 1184 31906 1193
rect 31850 1119 31906 1128
rect 29552 264 29604 270
rect 29552 206 29604 212
rect 26606 0 26662 40
rect 26790 0 26846 56
rect 26974 0 27030 56
rect 27158 0 27214 56
rect 27342 0 27398 56
rect 27526 0 27582 56
rect 27710 0 27766 56
rect 27894 54 28028 56
rect 27894 0 27950 54
rect 28078 0 28134 56
rect 28262 0 28318 56
rect 28446 0 28502 56
rect 28630 0 28686 56
<< via2 >>
rect 1306 9560 1362 9616
rect 846 4664 902 4720
rect 2778 8744 2834 8800
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 9176 8730 9232 8732
rect 9256 8730 9312 8732
rect 9016 8678 9062 8730
rect 9062 8678 9072 8730
rect 9096 8678 9126 8730
rect 9126 8678 9138 8730
rect 9138 8678 9152 8730
rect 9176 8678 9190 8730
rect 9190 8678 9202 8730
rect 9202 8678 9232 8730
rect 9256 8678 9266 8730
rect 9266 8678 9312 8730
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 9176 8676 9232 8678
rect 9256 8676 9312 8678
rect 2778 8336 2834 8392
rect 1766 8200 1822 8256
rect 1306 4936 1362 4992
rect 1306 4528 1362 4584
rect 1214 4392 1270 4448
rect 1122 4120 1178 4176
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 2594 7928 2650 7984
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 9176 7642 9232 7644
rect 9256 7642 9312 7644
rect 9016 7590 9062 7642
rect 9062 7590 9072 7642
rect 9096 7590 9126 7642
rect 9126 7590 9138 7642
rect 9138 7590 9152 7642
rect 9176 7590 9190 7642
rect 9190 7590 9202 7642
rect 9202 7590 9232 7642
rect 9256 7590 9266 7642
rect 9266 7590 9312 7642
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 9176 7588 9232 7590
rect 9256 7588 9312 7590
rect 14738 9016 14794 9072
rect 13956 8186 14012 8188
rect 14036 8186 14092 8188
rect 14116 8186 14172 8188
rect 14196 8186 14252 8188
rect 13956 8134 14002 8186
rect 14002 8134 14012 8186
rect 14036 8134 14066 8186
rect 14066 8134 14078 8186
rect 14078 8134 14092 8186
rect 14116 8134 14130 8186
rect 14130 8134 14142 8186
rect 14142 8134 14172 8186
rect 14196 8134 14206 8186
rect 14206 8134 14252 8186
rect 13956 8132 14012 8134
rect 14036 8132 14092 8134
rect 14116 8132 14172 8134
rect 14196 8132 14252 8134
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 1766 6024 1822 6080
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 1766 5616 1822 5672
rect 2870 6568 2926 6624
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 9176 6554 9232 6556
rect 9256 6554 9312 6556
rect 9016 6502 9062 6554
rect 9062 6502 9072 6554
rect 9096 6502 9126 6554
rect 9126 6502 9138 6554
rect 9138 6502 9152 6554
rect 9176 6502 9190 6554
rect 9190 6502 9202 6554
rect 9202 6502 9232 6554
rect 9256 6502 9266 6554
rect 9266 6502 9312 6554
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 9176 6500 9232 6502
rect 9256 6500 9312 6502
rect 2870 6160 2926 6216
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 13956 7098 14012 7100
rect 14036 7098 14092 7100
rect 14116 7098 14172 7100
rect 14196 7098 14252 7100
rect 13956 7046 14002 7098
rect 14002 7046 14012 7098
rect 14036 7046 14066 7098
rect 14066 7046 14078 7098
rect 14078 7046 14092 7098
rect 14116 7046 14130 7098
rect 14130 7046 14142 7098
rect 14142 7046 14172 7098
rect 14196 7046 14206 7098
rect 14206 7046 14252 7098
rect 13956 7044 14012 7046
rect 14036 7044 14092 7046
rect 14116 7044 14172 7046
rect 14196 7044 14252 7046
rect 13956 6010 14012 6012
rect 14036 6010 14092 6012
rect 14116 6010 14172 6012
rect 14196 6010 14252 6012
rect 13956 5958 14002 6010
rect 14002 5958 14012 6010
rect 14036 5958 14066 6010
rect 14066 5958 14078 6010
rect 14078 5958 14092 6010
rect 14116 5958 14130 6010
rect 14130 5958 14142 6010
rect 14142 5958 14172 6010
rect 14196 5958 14206 6010
rect 14206 5958 14252 6010
rect 13956 5956 14012 5958
rect 14036 5956 14092 5958
rect 14116 5956 14172 5958
rect 14196 5956 14252 5958
rect 2778 5480 2834 5536
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 9176 5466 9232 5468
rect 9256 5466 9312 5468
rect 9016 5414 9062 5466
rect 9062 5414 9072 5466
rect 9096 5414 9126 5466
rect 9126 5414 9138 5466
rect 9138 5414 9152 5466
rect 9176 5414 9190 5466
rect 9190 5414 9202 5466
rect 9202 5414 9232 5466
rect 9256 5414 9266 5466
rect 9266 5414 9312 5466
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 9176 5412 9232 5414
rect 9256 5412 9312 5414
rect 2686 5208 2742 5264
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 1674 3848 1730 3904
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 2502 3440 2558 3496
rect 1306 2760 1362 2816
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 2870 3304 2926 3360
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 2870 2896 2926 2952
rect 2870 2216 2926 2272
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 2870 1808 2926 1864
rect 4526 1264 4582 1320
rect 4894 40 4950 96
rect 7470 1264 7526 1320
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 7654 40 7710 96
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 9176 4378 9232 4380
rect 9256 4378 9312 4380
rect 9016 4326 9062 4378
rect 9062 4326 9072 4378
rect 9096 4326 9126 4378
rect 9126 4326 9138 4378
rect 9138 4326 9152 4378
rect 9176 4326 9190 4378
rect 9190 4326 9202 4378
rect 9202 4326 9232 4378
rect 9256 4326 9266 4378
rect 9266 4326 9312 4378
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 9176 4324 9232 4326
rect 9256 4324 9312 4326
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 9176 3290 9232 3292
rect 9256 3290 9312 3292
rect 9016 3238 9062 3290
rect 9062 3238 9072 3290
rect 9096 3238 9126 3290
rect 9126 3238 9138 3290
rect 9138 3238 9152 3290
rect 9176 3238 9190 3290
rect 9190 3238 9202 3290
rect 9202 3238 9232 3290
rect 9256 3238 9266 3290
rect 9266 3238 9312 3290
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 9176 3236 9232 3238
rect 9256 3236 9312 3238
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 9176 2202 9232 2204
rect 9256 2202 9312 2204
rect 9016 2150 9062 2202
rect 9062 2150 9072 2202
rect 9096 2150 9126 2202
rect 9126 2150 9138 2202
rect 9138 2150 9152 2202
rect 9176 2150 9190 2202
rect 9190 2150 9202 2202
rect 9202 2150 9232 2202
rect 9256 2150 9266 2202
rect 9266 2150 9312 2202
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 9176 2148 9232 2150
rect 9256 2148 9312 2150
rect 9862 2080 9918 2136
rect 11058 5072 11114 5128
rect 11610 4664 11666 4720
rect 12438 2352 12494 2408
rect 15016 8730 15072 8732
rect 15096 8730 15152 8732
rect 15176 8730 15232 8732
rect 15256 8730 15312 8732
rect 15016 8678 15062 8730
rect 15062 8678 15072 8730
rect 15096 8678 15126 8730
rect 15126 8678 15138 8730
rect 15138 8678 15152 8730
rect 15176 8678 15190 8730
rect 15190 8678 15202 8730
rect 15202 8678 15232 8730
rect 15256 8678 15266 8730
rect 15266 8678 15312 8730
rect 15016 8676 15072 8678
rect 15096 8676 15152 8678
rect 15176 8676 15232 8678
rect 15256 8676 15312 8678
rect 16946 9288 17002 9344
rect 15016 7642 15072 7644
rect 15096 7642 15152 7644
rect 15176 7642 15232 7644
rect 15256 7642 15312 7644
rect 15016 7590 15062 7642
rect 15062 7590 15072 7642
rect 15096 7590 15126 7642
rect 15126 7590 15138 7642
rect 15138 7590 15152 7642
rect 15176 7590 15190 7642
rect 15190 7590 15202 7642
rect 15202 7590 15232 7642
rect 15256 7590 15266 7642
rect 15266 7590 15312 7642
rect 15016 7588 15072 7590
rect 15096 7588 15152 7590
rect 15176 7588 15232 7590
rect 15256 7588 15312 7590
rect 15474 7384 15530 7440
rect 13956 4922 14012 4924
rect 14036 4922 14092 4924
rect 14116 4922 14172 4924
rect 14196 4922 14252 4924
rect 13956 4870 14002 4922
rect 14002 4870 14012 4922
rect 14036 4870 14066 4922
rect 14066 4870 14078 4922
rect 14078 4870 14092 4922
rect 14116 4870 14130 4922
rect 14130 4870 14142 4922
rect 14142 4870 14172 4922
rect 14196 4870 14206 4922
rect 14206 4870 14252 4922
rect 13956 4868 14012 4870
rect 14036 4868 14092 4870
rect 14116 4868 14172 4870
rect 14196 4868 14252 4870
rect 13956 3834 14012 3836
rect 14036 3834 14092 3836
rect 14116 3834 14172 3836
rect 14196 3834 14252 3836
rect 13956 3782 14002 3834
rect 14002 3782 14012 3834
rect 14036 3782 14066 3834
rect 14066 3782 14078 3834
rect 14078 3782 14092 3834
rect 14116 3782 14130 3834
rect 14130 3782 14142 3834
rect 14142 3782 14172 3834
rect 14196 3782 14206 3834
rect 14206 3782 14252 3834
rect 13956 3780 14012 3782
rect 14036 3780 14092 3782
rect 14116 3780 14172 3782
rect 14196 3780 14252 3782
rect 14462 3848 14518 3904
rect 13956 2746 14012 2748
rect 14036 2746 14092 2748
rect 14116 2746 14172 2748
rect 14196 2746 14252 2748
rect 13956 2694 14002 2746
rect 14002 2694 14012 2746
rect 14036 2694 14066 2746
rect 14066 2694 14078 2746
rect 14078 2694 14092 2746
rect 14116 2694 14130 2746
rect 14130 2694 14142 2746
rect 14142 2694 14172 2746
rect 14196 2694 14206 2746
rect 14206 2694 14252 2746
rect 13956 2692 14012 2694
rect 14036 2692 14092 2694
rect 14116 2692 14172 2694
rect 14196 2692 14252 2694
rect 13818 2080 13874 2136
rect 13726 584 13782 640
rect 13542 448 13598 504
rect 13358 312 13414 368
rect 13910 176 13966 232
rect 14738 3984 14794 4040
rect 14830 2760 14886 2816
rect 15016 6554 15072 6556
rect 15096 6554 15152 6556
rect 15176 6554 15232 6556
rect 15256 6554 15312 6556
rect 15016 6502 15062 6554
rect 15062 6502 15072 6554
rect 15096 6502 15126 6554
rect 15126 6502 15138 6554
rect 15138 6502 15152 6554
rect 15176 6502 15190 6554
rect 15190 6502 15202 6554
rect 15202 6502 15232 6554
rect 15256 6502 15266 6554
rect 15266 6502 15312 6554
rect 15016 6500 15072 6502
rect 15096 6500 15152 6502
rect 15176 6500 15232 6502
rect 15256 6500 15312 6502
rect 15106 6332 15108 6352
rect 15108 6332 15160 6352
rect 15160 6332 15162 6352
rect 15106 6296 15162 6332
rect 15016 5466 15072 5468
rect 15096 5466 15152 5468
rect 15176 5466 15232 5468
rect 15256 5466 15312 5468
rect 15016 5414 15062 5466
rect 15062 5414 15072 5466
rect 15096 5414 15126 5466
rect 15126 5414 15138 5466
rect 15138 5414 15152 5466
rect 15176 5414 15190 5466
rect 15190 5414 15202 5466
rect 15202 5414 15232 5466
rect 15256 5414 15266 5466
rect 15266 5414 15312 5466
rect 15016 5412 15072 5414
rect 15096 5412 15152 5414
rect 15176 5412 15232 5414
rect 15256 5412 15312 5414
rect 16486 7248 16542 7304
rect 15750 6840 15806 6896
rect 15658 5072 15714 5128
rect 15016 4378 15072 4380
rect 15096 4378 15152 4380
rect 15176 4378 15232 4380
rect 15256 4378 15312 4380
rect 15016 4326 15062 4378
rect 15062 4326 15072 4378
rect 15096 4326 15126 4378
rect 15126 4326 15138 4378
rect 15138 4326 15152 4378
rect 15176 4326 15190 4378
rect 15190 4326 15202 4378
rect 15202 4326 15232 4378
rect 15256 4326 15266 4378
rect 15266 4326 15312 4378
rect 15016 4324 15072 4326
rect 15096 4324 15152 4326
rect 15176 4324 15232 4326
rect 15256 4324 15312 4326
rect 15016 3290 15072 3292
rect 15096 3290 15152 3292
rect 15176 3290 15232 3292
rect 15256 3290 15312 3292
rect 15016 3238 15062 3290
rect 15062 3238 15072 3290
rect 15096 3238 15126 3290
rect 15126 3238 15138 3290
rect 15138 3238 15152 3290
rect 15176 3238 15190 3290
rect 15190 3238 15202 3290
rect 15202 3238 15232 3290
rect 15256 3238 15266 3290
rect 15266 3238 15312 3290
rect 15016 3236 15072 3238
rect 15096 3236 15152 3238
rect 15176 3236 15232 3238
rect 15256 3236 15312 3238
rect 16210 6160 16266 6216
rect 15934 5208 15990 5264
rect 16394 5616 16450 5672
rect 15016 2202 15072 2204
rect 15096 2202 15152 2204
rect 15176 2202 15232 2204
rect 15256 2202 15312 2204
rect 15016 2150 15062 2202
rect 15062 2150 15072 2202
rect 15096 2150 15126 2202
rect 15126 2150 15138 2202
rect 15138 2150 15152 2202
rect 15176 2150 15190 2202
rect 15190 2150 15202 2202
rect 15202 2150 15232 2202
rect 15256 2150 15266 2202
rect 15266 2150 15312 2202
rect 15016 2148 15072 2150
rect 15096 2148 15152 2150
rect 15176 2148 15232 2150
rect 15256 2148 15312 2150
rect 16026 2760 16082 2816
rect 17038 8472 17094 8528
rect 17498 8336 17554 8392
rect 18970 7792 19026 7848
rect 17130 4528 17186 4584
rect 16762 3440 16818 3496
rect 16762 1672 16818 1728
rect 17498 1808 17554 1864
rect 17682 1128 17738 1184
rect 21016 8730 21072 8732
rect 21096 8730 21152 8732
rect 21176 8730 21232 8732
rect 21256 8730 21312 8732
rect 21016 8678 21062 8730
rect 21062 8678 21072 8730
rect 21096 8678 21126 8730
rect 21126 8678 21138 8730
rect 21138 8678 21152 8730
rect 21176 8678 21190 8730
rect 21190 8678 21202 8730
rect 21202 8678 21232 8730
rect 21256 8678 21266 8730
rect 21266 8678 21312 8730
rect 21016 8676 21072 8678
rect 21096 8676 21152 8678
rect 21176 8676 21232 8678
rect 21256 8676 21312 8678
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 20196 8186 20252 8188
rect 19956 8134 20002 8186
rect 20002 8134 20012 8186
rect 20036 8134 20066 8186
rect 20066 8134 20078 8186
rect 20078 8134 20092 8186
rect 20116 8134 20130 8186
rect 20130 8134 20142 8186
rect 20142 8134 20172 8186
rect 20196 8134 20206 8186
rect 20206 8134 20252 8186
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 20196 8132 20252 8134
rect 21016 7642 21072 7644
rect 21096 7642 21152 7644
rect 21176 7642 21232 7644
rect 21256 7642 21312 7644
rect 21016 7590 21062 7642
rect 21062 7590 21072 7642
rect 21096 7590 21126 7642
rect 21126 7590 21138 7642
rect 21138 7590 21152 7642
rect 21176 7590 21190 7642
rect 21190 7590 21202 7642
rect 21202 7590 21232 7642
rect 21256 7590 21266 7642
rect 21266 7590 21312 7642
rect 21016 7588 21072 7590
rect 21096 7588 21152 7590
rect 21176 7588 21232 7590
rect 21256 7588 21312 7590
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 20196 7098 20252 7100
rect 19956 7046 20002 7098
rect 20002 7046 20012 7098
rect 20036 7046 20066 7098
rect 20066 7046 20078 7098
rect 20078 7046 20092 7098
rect 20116 7046 20130 7098
rect 20130 7046 20142 7098
rect 20142 7046 20172 7098
rect 20196 7046 20206 7098
rect 20206 7046 20252 7098
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 20196 7044 20252 7046
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 20196 6010 20252 6012
rect 19956 5958 20002 6010
rect 20002 5958 20012 6010
rect 20036 5958 20066 6010
rect 20066 5958 20078 6010
rect 20078 5958 20092 6010
rect 20116 5958 20130 6010
rect 20130 5958 20142 6010
rect 20142 5958 20172 6010
rect 20196 5958 20206 6010
rect 20206 5958 20252 6010
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 20196 5956 20252 5958
rect 21016 6554 21072 6556
rect 21096 6554 21152 6556
rect 21176 6554 21232 6556
rect 21256 6554 21312 6556
rect 21016 6502 21062 6554
rect 21062 6502 21072 6554
rect 21096 6502 21126 6554
rect 21126 6502 21138 6554
rect 21138 6502 21152 6554
rect 21176 6502 21190 6554
rect 21190 6502 21202 6554
rect 21202 6502 21232 6554
rect 21256 6502 21266 6554
rect 21266 6502 21312 6554
rect 21016 6500 21072 6502
rect 21096 6500 21152 6502
rect 21176 6500 21232 6502
rect 21256 6500 21312 6502
rect 21016 5466 21072 5468
rect 21096 5466 21152 5468
rect 21176 5466 21232 5468
rect 21256 5466 21312 5468
rect 21016 5414 21062 5466
rect 21062 5414 21072 5466
rect 21096 5414 21126 5466
rect 21126 5414 21138 5466
rect 21138 5414 21152 5466
rect 21176 5414 21190 5466
rect 21190 5414 21202 5466
rect 21202 5414 21232 5466
rect 21256 5414 21266 5466
rect 21266 5414 21312 5466
rect 21016 5412 21072 5414
rect 21096 5412 21152 5414
rect 21176 5412 21232 5414
rect 21256 5412 21312 5414
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 20196 4922 20252 4924
rect 19956 4870 20002 4922
rect 20002 4870 20012 4922
rect 20036 4870 20066 4922
rect 20066 4870 20078 4922
rect 20078 4870 20092 4922
rect 20116 4870 20130 4922
rect 20130 4870 20142 4922
rect 20142 4870 20172 4922
rect 20196 4870 20206 4922
rect 20206 4870 20252 4922
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 20196 4868 20252 4870
rect 20810 4664 20866 4720
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 20196 3834 20252 3836
rect 19956 3782 20002 3834
rect 20002 3782 20012 3834
rect 20036 3782 20066 3834
rect 20066 3782 20078 3834
rect 20078 3782 20092 3834
rect 20116 3782 20130 3834
rect 20130 3782 20142 3834
rect 20142 3782 20172 3834
rect 20196 3782 20206 3834
rect 20206 3782 20252 3834
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 20196 3780 20252 3782
rect 20718 3596 20774 3632
rect 20718 3576 20720 3596
rect 20720 3576 20772 3596
rect 20772 3576 20774 3596
rect 19430 1400 19486 1456
rect 19706 1808 19762 1864
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 20196 2746 20252 2748
rect 19956 2694 20002 2746
rect 20002 2694 20012 2746
rect 20036 2694 20066 2746
rect 20066 2694 20078 2746
rect 20078 2694 20092 2746
rect 20116 2694 20130 2746
rect 20130 2694 20142 2746
rect 20142 2694 20172 2746
rect 20196 2694 20206 2746
rect 20206 2694 20252 2746
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 20196 2692 20252 2694
rect 21016 4378 21072 4380
rect 21096 4378 21152 4380
rect 21176 4378 21232 4380
rect 21256 4378 21312 4380
rect 21016 4326 21062 4378
rect 21062 4326 21072 4378
rect 21096 4326 21126 4378
rect 21126 4326 21138 4378
rect 21138 4326 21152 4378
rect 21176 4326 21190 4378
rect 21190 4326 21202 4378
rect 21202 4326 21232 4378
rect 21256 4326 21266 4378
rect 21266 4326 21312 4378
rect 21016 4324 21072 4326
rect 21096 4324 21152 4326
rect 21176 4324 21232 4326
rect 21256 4324 21312 4326
rect 21016 3290 21072 3292
rect 21096 3290 21152 3292
rect 21176 3290 21232 3292
rect 21256 3290 21312 3292
rect 21016 3238 21062 3290
rect 21062 3238 21072 3290
rect 21096 3238 21126 3290
rect 21126 3238 21138 3290
rect 21138 3238 21152 3290
rect 21176 3238 21190 3290
rect 21190 3238 21202 3290
rect 21202 3238 21232 3290
rect 21256 3238 21266 3290
rect 21266 3238 21312 3290
rect 21016 3236 21072 3238
rect 21096 3236 21152 3238
rect 21176 3236 21232 3238
rect 21256 3236 21312 3238
rect 21638 3340 21640 3360
rect 21640 3340 21692 3360
rect 21692 3340 21694 3360
rect 21638 3304 21694 3340
rect 21016 2202 21072 2204
rect 21096 2202 21152 2204
rect 21176 2202 21232 2204
rect 21256 2202 21312 2204
rect 21016 2150 21062 2202
rect 21062 2150 21072 2202
rect 21096 2150 21126 2202
rect 21126 2150 21138 2202
rect 21138 2150 21152 2202
rect 21176 2150 21190 2202
rect 21190 2150 21202 2202
rect 21202 2150 21232 2202
rect 21256 2150 21266 2202
rect 21266 2150 21312 2202
rect 21016 2148 21072 2150
rect 21096 2148 21152 2150
rect 21176 2148 21232 2150
rect 21256 2148 21312 2150
rect 22282 5752 22338 5808
rect 22190 3340 22192 3360
rect 22192 3340 22244 3360
rect 22244 3340 22246 3360
rect 21914 1944 21970 2000
rect 22190 3304 22246 3340
rect 24858 5788 24860 5808
rect 24860 5788 24912 5808
rect 24912 5788 24914 5808
rect 24858 5752 24914 5788
rect 23018 2624 23074 2680
rect 23570 3032 23626 3088
rect 23386 2488 23442 2544
rect 24122 3440 24178 3496
rect 23938 2488 23994 2544
rect 24582 3032 24638 3088
rect 24766 3612 24768 3632
rect 24768 3612 24820 3632
rect 24820 3612 24822 3632
rect 24766 3576 24822 3612
rect 24858 2896 24914 2952
rect 25318 1808 25374 1864
rect 25134 40 25190 96
rect 25502 2624 25558 2680
rect 25594 1264 25650 1320
rect 25410 40 25466 96
rect 27016 8730 27072 8732
rect 27096 8730 27152 8732
rect 27176 8730 27232 8732
rect 27256 8730 27312 8732
rect 27016 8678 27062 8730
rect 27062 8678 27072 8730
rect 27096 8678 27126 8730
rect 27126 8678 27138 8730
rect 27138 8678 27152 8730
rect 27176 8678 27190 8730
rect 27190 8678 27202 8730
rect 27202 8678 27232 8730
rect 27256 8678 27266 8730
rect 27266 8678 27312 8730
rect 27016 8676 27072 8678
rect 27096 8676 27152 8678
rect 27176 8676 27232 8678
rect 27256 8676 27312 8678
rect 25956 8186 26012 8188
rect 26036 8186 26092 8188
rect 26116 8186 26172 8188
rect 26196 8186 26252 8188
rect 25956 8134 26002 8186
rect 26002 8134 26012 8186
rect 26036 8134 26066 8186
rect 26066 8134 26078 8186
rect 26078 8134 26092 8186
rect 26116 8134 26130 8186
rect 26130 8134 26142 8186
rect 26142 8134 26172 8186
rect 26196 8134 26206 8186
rect 26206 8134 26252 8186
rect 25956 8132 26012 8134
rect 26036 8132 26092 8134
rect 26116 8132 26172 8134
rect 26196 8132 26252 8134
rect 27016 7642 27072 7644
rect 27096 7642 27152 7644
rect 27176 7642 27232 7644
rect 27256 7642 27312 7644
rect 27016 7590 27062 7642
rect 27062 7590 27072 7642
rect 27096 7590 27126 7642
rect 27126 7590 27138 7642
rect 27138 7590 27152 7642
rect 27176 7590 27190 7642
rect 27190 7590 27202 7642
rect 27202 7590 27232 7642
rect 27256 7590 27266 7642
rect 27266 7590 27312 7642
rect 27016 7588 27072 7590
rect 27096 7588 27152 7590
rect 27176 7588 27232 7590
rect 27256 7588 27312 7590
rect 31114 9288 31170 9344
rect 25956 7098 26012 7100
rect 26036 7098 26092 7100
rect 26116 7098 26172 7100
rect 26196 7098 26252 7100
rect 25956 7046 26002 7098
rect 26002 7046 26012 7098
rect 26036 7046 26066 7098
rect 26066 7046 26078 7098
rect 26078 7046 26092 7098
rect 26116 7046 26130 7098
rect 26130 7046 26142 7098
rect 26142 7046 26172 7098
rect 26196 7046 26206 7098
rect 26206 7046 26252 7098
rect 25956 7044 26012 7046
rect 26036 7044 26092 7046
rect 26116 7044 26172 7046
rect 26196 7044 26252 7046
rect 25956 6010 26012 6012
rect 26036 6010 26092 6012
rect 26116 6010 26172 6012
rect 26196 6010 26252 6012
rect 25956 5958 26002 6010
rect 26002 5958 26012 6010
rect 26036 5958 26066 6010
rect 26066 5958 26078 6010
rect 26078 5958 26092 6010
rect 26116 5958 26130 6010
rect 26130 5958 26142 6010
rect 26142 5958 26172 6010
rect 26196 5958 26206 6010
rect 26206 5958 26252 6010
rect 25956 5956 26012 5958
rect 26036 5956 26092 5958
rect 26116 5956 26172 5958
rect 26196 5956 26252 5958
rect 25956 4922 26012 4924
rect 26036 4922 26092 4924
rect 26116 4922 26172 4924
rect 26196 4922 26252 4924
rect 25956 4870 26002 4922
rect 26002 4870 26012 4922
rect 26036 4870 26066 4922
rect 26066 4870 26078 4922
rect 26078 4870 26092 4922
rect 26116 4870 26130 4922
rect 26130 4870 26142 4922
rect 26142 4870 26172 4922
rect 26196 4870 26206 4922
rect 26206 4870 26252 4922
rect 25956 4868 26012 4870
rect 26036 4868 26092 4870
rect 26116 4868 26172 4870
rect 26196 4868 26252 4870
rect 25956 3834 26012 3836
rect 26036 3834 26092 3836
rect 26116 3834 26172 3836
rect 26196 3834 26252 3836
rect 25956 3782 26002 3834
rect 26002 3782 26012 3834
rect 26036 3782 26066 3834
rect 26066 3782 26078 3834
rect 26078 3782 26092 3834
rect 26116 3782 26130 3834
rect 26130 3782 26142 3834
rect 26142 3782 26172 3834
rect 26196 3782 26206 3834
rect 26206 3782 26252 3834
rect 25956 3780 26012 3782
rect 26036 3780 26092 3782
rect 26116 3780 26172 3782
rect 26196 3780 26252 3782
rect 26330 3712 26386 3768
rect 25956 2746 26012 2748
rect 26036 2746 26092 2748
rect 26116 2746 26172 2748
rect 26196 2746 26252 2748
rect 25956 2694 26002 2746
rect 26002 2694 26012 2746
rect 26036 2694 26066 2746
rect 26066 2694 26078 2746
rect 26078 2694 26092 2746
rect 26116 2694 26130 2746
rect 26130 2694 26142 2746
rect 26142 2694 26172 2746
rect 26196 2694 26206 2746
rect 26206 2694 26252 2746
rect 25956 2692 26012 2694
rect 26036 2692 26092 2694
rect 26116 2692 26172 2694
rect 26196 2692 26252 2694
rect 25778 2488 25834 2544
rect 26054 2488 26110 2544
rect 26698 5208 26754 5264
rect 27016 6554 27072 6556
rect 27096 6554 27152 6556
rect 27176 6554 27232 6556
rect 27256 6554 27312 6556
rect 27016 6502 27062 6554
rect 27062 6502 27072 6554
rect 27096 6502 27126 6554
rect 27126 6502 27138 6554
rect 27138 6502 27152 6554
rect 27176 6502 27190 6554
rect 27190 6502 27202 6554
rect 27202 6502 27232 6554
rect 27256 6502 27266 6554
rect 27266 6502 27312 6554
rect 27016 6500 27072 6502
rect 27096 6500 27152 6502
rect 27176 6500 27232 6502
rect 27256 6500 27312 6502
rect 27016 5466 27072 5468
rect 27096 5466 27152 5468
rect 27176 5466 27232 5468
rect 27256 5466 27312 5468
rect 27016 5414 27062 5466
rect 27062 5414 27072 5466
rect 27096 5414 27126 5466
rect 27126 5414 27138 5466
rect 27138 5414 27152 5466
rect 27176 5414 27190 5466
rect 27190 5414 27202 5466
rect 27202 5414 27232 5466
rect 27256 5414 27266 5466
rect 27266 5414 27312 5466
rect 27016 5412 27072 5414
rect 27096 5412 27152 5414
rect 27176 5412 27232 5414
rect 27256 5412 27312 5414
rect 27016 4378 27072 4380
rect 27096 4378 27152 4380
rect 27176 4378 27232 4380
rect 27256 4378 27312 4380
rect 27016 4326 27062 4378
rect 27062 4326 27072 4378
rect 27096 4326 27126 4378
rect 27126 4326 27138 4378
rect 27138 4326 27152 4378
rect 27176 4326 27190 4378
rect 27190 4326 27202 4378
rect 27202 4326 27232 4378
rect 27256 4326 27266 4378
rect 27266 4326 27312 4378
rect 27016 4324 27072 4326
rect 27096 4324 27152 4326
rect 27176 4324 27232 4326
rect 27256 4324 27312 4326
rect 27526 4120 27582 4176
rect 27016 3290 27072 3292
rect 27096 3290 27152 3292
rect 27176 3290 27232 3292
rect 27256 3290 27312 3292
rect 27016 3238 27062 3290
rect 27062 3238 27072 3290
rect 27096 3238 27126 3290
rect 27126 3238 27138 3290
rect 27138 3238 27152 3290
rect 27176 3238 27190 3290
rect 27190 3238 27202 3290
rect 27202 3238 27232 3290
rect 27256 3238 27266 3290
rect 27266 3238 27312 3290
rect 27016 3236 27072 3238
rect 27096 3236 27152 3238
rect 27176 3236 27232 3238
rect 27256 3236 27312 3238
rect 26882 2352 26938 2408
rect 26606 40 26662 96
rect 27016 2202 27072 2204
rect 27096 2202 27152 2204
rect 27176 2202 27232 2204
rect 27256 2202 27312 2204
rect 27016 2150 27062 2202
rect 27062 2150 27072 2202
rect 27096 2150 27126 2202
rect 27126 2150 27138 2202
rect 27138 2150 27152 2202
rect 27176 2150 27190 2202
rect 27190 2150 27202 2202
rect 27202 2150 27232 2202
rect 27256 2150 27266 2202
rect 27266 2150 27312 2202
rect 27016 2148 27072 2150
rect 27096 2148 27152 2150
rect 27176 2148 27232 2150
rect 27256 2148 27312 2150
rect 26974 1264 27030 1320
rect 26882 312 26938 368
rect 27526 1400 27582 1456
rect 27894 4120 27950 4176
rect 27802 2896 27858 2952
rect 28446 4664 28502 4720
rect 28262 4564 28264 4584
rect 28264 4564 28316 4584
rect 28316 4564 28318 4584
rect 28262 4528 28318 4564
rect 28446 4020 28448 4040
rect 28448 4020 28500 4040
rect 28500 4020 28502 4040
rect 28446 3984 28502 4020
rect 28262 3440 28318 3496
rect 28446 3068 28448 3088
rect 28448 3068 28500 3088
rect 28500 3068 28502 3088
rect 28446 3032 28502 3068
rect 30378 3596 30434 3632
rect 30378 3576 30380 3596
rect 30380 3576 30432 3596
rect 30432 3576 30434 3596
rect 31390 9560 31446 9616
rect 31758 9016 31814 9072
rect 33414 8744 33470 8800
rect 33016 8730 33072 8732
rect 33096 8730 33152 8732
rect 33176 8730 33232 8732
rect 33256 8730 33312 8732
rect 33016 8678 33062 8730
rect 33062 8678 33072 8730
rect 33096 8678 33126 8730
rect 33126 8678 33138 8730
rect 33138 8678 33152 8730
rect 33176 8678 33190 8730
rect 33190 8678 33202 8730
rect 33202 8678 33232 8730
rect 33256 8678 33266 8730
rect 33266 8678 33312 8730
rect 33016 8676 33072 8678
rect 33096 8676 33152 8678
rect 33176 8676 33232 8678
rect 33256 8676 33312 8678
rect 32310 8472 32366 8528
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 33046 8200 33102 8256
rect 32494 7928 32550 7984
rect 33016 7642 33072 7644
rect 33096 7642 33152 7644
rect 33176 7642 33232 7644
rect 33256 7642 33312 7644
rect 33016 7590 33062 7642
rect 33062 7590 33072 7642
rect 33096 7590 33126 7642
rect 33126 7590 33138 7642
rect 33138 7590 33152 7642
rect 33176 7590 33190 7642
rect 33190 7590 33202 7642
rect 33202 7590 33232 7642
rect 33256 7590 33266 7642
rect 33266 7590 33312 7642
rect 33016 7588 33072 7590
rect 33096 7588 33152 7590
rect 33176 7588 33232 7590
rect 33256 7588 33312 7590
rect 33598 7692 33600 7712
rect 33600 7692 33652 7712
rect 33652 7692 33654 7712
rect 33598 7656 33654 7692
rect 32494 7384 32550 7440
rect 32862 7148 32864 7168
rect 32864 7148 32916 7168
rect 32916 7148 32918 7168
rect 32862 7112 32918 7148
rect 32862 6840 32918 6896
rect 33414 6568 33470 6624
rect 33016 6554 33072 6556
rect 33096 6554 33152 6556
rect 33176 6554 33232 6556
rect 33256 6554 33312 6556
rect 33016 6502 33062 6554
rect 33062 6502 33072 6554
rect 33096 6502 33126 6554
rect 33126 6502 33138 6554
rect 33138 6502 33152 6554
rect 33176 6502 33190 6554
rect 33190 6502 33202 6554
rect 33202 6502 33232 6554
rect 33256 6502 33266 6554
rect 33266 6502 33312 6554
rect 33016 6500 33072 6502
rect 33096 6500 33152 6502
rect 33176 6500 33232 6502
rect 33256 6500 33312 6502
rect 32862 6296 32918 6352
rect 32494 6060 32496 6080
rect 32496 6060 32548 6080
rect 32548 6060 32550 6080
rect 32494 6024 32550 6060
rect 32862 5788 32864 5808
rect 32864 5788 32916 5808
rect 32916 5788 32918 5808
rect 32862 5752 32918 5788
rect 33414 5516 33416 5536
rect 33416 5516 33468 5536
rect 33468 5516 33470 5536
rect 33414 5480 33470 5516
rect 33016 5466 33072 5468
rect 33096 5466 33152 5468
rect 33176 5466 33232 5468
rect 33256 5466 33312 5468
rect 33016 5414 33062 5466
rect 33062 5414 33072 5466
rect 33096 5414 33126 5466
rect 33126 5414 33138 5466
rect 33138 5414 33152 5466
rect 33176 5414 33190 5466
rect 33190 5414 33202 5466
rect 33202 5414 33232 5466
rect 33256 5414 33266 5466
rect 33266 5414 33312 5466
rect 33016 5412 33072 5414
rect 33096 5412 33152 5414
rect 33176 5412 33232 5414
rect 33256 5412 33312 5414
rect 32862 5208 32918 5264
rect 32494 4972 32496 4992
rect 32496 4972 32548 4992
rect 32548 4972 32550 4992
rect 32494 4936 32550 4972
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 32862 4700 32864 4720
rect 32864 4700 32916 4720
rect 32916 4700 32918 4720
rect 32862 4664 32918 4700
rect 33414 4428 33416 4448
rect 33416 4428 33468 4448
rect 33468 4428 33470 4448
rect 33414 4392 33470 4428
rect 33016 4378 33072 4380
rect 33096 4378 33152 4380
rect 33176 4378 33232 4380
rect 33256 4378 33312 4380
rect 33016 4326 33062 4378
rect 33062 4326 33072 4378
rect 33096 4326 33126 4378
rect 33126 4326 33138 4378
rect 33138 4326 33152 4378
rect 33176 4326 33190 4378
rect 33190 4326 33202 4378
rect 33202 4326 33232 4378
rect 33256 4326 33266 4378
rect 33266 4326 33312 4378
rect 33016 4324 33072 4326
rect 33096 4324 33152 4326
rect 33176 4324 33232 4326
rect 33256 4324 33312 4326
rect 32862 4120 32918 4176
rect 32494 3884 32496 3904
rect 32496 3884 32548 3904
rect 32548 3884 32550 3904
rect 32494 3848 32550 3884
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 31666 3712 31722 3768
rect 32862 3612 32864 3632
rect 32864 3612 32916 3632
rect 32916 3612 32918 3632
rect 32862 3576 32918 3612
rect 33414 3340 33416 3360
rect 33416 3340 33468 3360
rect 33468 3340 33470 3360
rect 33414 3304 33470 3340
rect 33016 3290 33072 3292
rect 33096 3290 33152 3292
rect 33176 3290 33232 3292
rect 33256 3290 33312 3292
rect 33016 3238 33062 3290
rect 33062 3238 33072 3290
rect 33096 3238 33126 3290
rect 33126 3238 33138 3290
rect 33138 3238 33152 3290
rect 33176 3238 33190 3290
rect 33190 3238 33202 3290
rect 33202 3238 33232 3290
rect 33256 3238 33266 3290
rect 33266 3238 33312 3290
rect 33016 3236 33072 3238
rect 33096 3236 33152 3238
rect 33176 3236 33232 3238
rect 33256 3236 33312 3238
rect 32862 3032 32918 3088
rect 32494 2796 32496 2816
rect 32496 2796 32548 2816
rect 32548 2796 32550 2816
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 31114 1944 31170 2000
rect 30470 1400 30526 1456
rect 31482 1400 31538 1456
rect 32494 2760 32550 2796
rect 32862 2524 32864 2544
rect 32864 2524 32916 2544
rect 32916 2524 32918 2544
rect 32862 2488 32918 2524
rect 33414 2252 33416 2272
rect 33416 2252 33468 2272
rect 33468 2252 33470 2272
rect 33414 2216 33470 2252
rect 33016 2202 33072 2204
rect 33096 2202 33152 2204
rect 33176 2202 33232 2204
rect 33256 2202 33312 2204
rect 33016 2150 33062 2202
rect 33062 2150 33072 2202
rect 33096 2150 33126 2202
rect 33126 2150 33138 2202
rect 33138 2150 33152 2202
rect 33176 2150 33190 2202
rect 33190 2150 33202 2202
rect 33202 2150 33232 2202
rect 33256 2150 33266 2202
rect 33266 2150 33312 2202
rect 33016 2148 33072 2150
rect 33096 2148 33152 2150
rect 33176 2148 33232 2150
rect 33256 2148 33312 2150
rect 32402 1672 32458 1728
rect 31850 1128 31906 1184
<< metal3 >>
rect 0 9618 120 9648
rect 1301 9618 1367 9621
rect 0 9616 1367 9618
rect 0 9560 1306 9616
rect 1362 9560 1367 9616
rect 0 9558 1367 9560
rect 0 9528 120 9558
rect 1301 9555 1367 9558
rect 31385 9618 31451 9621
rect 34288 9618 34408 9648
rect 31385 9616 34408 9618
rect 31385 9560 31390 9616
rect 31446 9560 34408 9616
rect 31385 9558 34408 9560
rect 31385 9555 31451 9558
rect 34288 9528 34408 9558
rect 0 9346 120 9376
rect 16941 9346 17007 9349
rect 0 9344 17007 9346
rect 0 9288 16946 9344
rect 17002 9288 17007 9344
rect 0 9286 17007 9288
rect 0 9256 120 9286
rect 16941 9283 17007 9286
rect 31109 9346 31175 9349
rect 34288 9346 34408 9376
rect 31109 9344 34408 9346
rect 31109 9288 31114 9344
rect 31170 9288 34408 9344
rect 31109 9286 34408 9288
rect 31109 9283 31175 9286
rect 34288 9256 34408 9286
rect 0 9074 120 9104
rect 14733 9074 14799 9077
rect 0 9072 14799 9074
rect 0 9016 14738 9072
rect 14794 9016 14799 9072
rect 0 9014 14799 9016
rect 0 8984 120 9014
rect 14733 9011 14799 9014
rect 31753 9074 31819 9077
rect 34288 9074 34408 9104
rect 31753 9072 34408 9074
rect 31753 9016 31758 9072
rect 31814 9016 34408 9072
rect 31753 9014 34408 9016
rect 31753 9011 31819 9014
rect 34288 8984 34408 9014
rect 0 8802 120 8832
rect 2773 8802 2839 8805
rect 0 8800 2839 8802
rect 0 8744 2778 8800
rect 2834 8744 2839 8800
rect 0 8742 2839 8744
rect 0 8712 120 8742
rect 2773 8739 2839 8742
rect 33409 8802 33475 8805
rect 34288 8802 34408 8832
rect 33409 8800 34408 8802
rect 33409 8744 33414 8800
rect 33470 8744 34408 8800
rect 33409 8742 34408 8744
rect 33409 8739 33475 8742
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 9006 8736 9322 8737
rect 9006 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9322 8736
rect 9006 8671 9322 8672
rect 15006 8736 15322 8737
rect 15006 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15322 8736
rect 15006 8671 15322 8672
rect 21006 8736 21322 8737
rect 21006 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21322 8736
rect 21006 8671 21322 8672
rect 27006 8736 27322 8737
rect 27006 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27322 8736
rect 27006 8671 27322 8672
rect 33006 8736 33322 8737
rect 33006 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33322 8736
rect 34288 8712 34408 8742
rect 33006 8671 33322 8672
rect 0 8530 120 8560
rect 17033 8530 17099 8533
rect 0 8528 17099 8530
rect 0 8472 17038 8528
rect 17094 8472 17099 8528
rect 0 8470 17099 8472
rect 0 8440 120 8470
rect 17033 8467 17099 8470
rect 32305 8530 32371 8533
rect 34288 8530 34408 8560
rect 32305 8528 34408 8530
rect 32305 8472 32310 8528
rect 32366 8472 34408 8528
rect 32305 8470 34408 8472
rect 32305 8467 32371 8470
rect 34288 8440 34408 8470
rect 2773 8394 2839 8397
rect 17493 8394 17559 8397
rect 2773 8392 17559 8394
rect 2773 8336 2778 8392
rect 2834 8336 17498 8392
rect 17554 8336 17559 8392
rect 2773 8334 17559 8336
rect 2773 8331 2839 8334
rect 17493 8331 17559 8334
rect 0 8258 120 8288
rect 1761 8258 1827 8261
rect 0 8256 1827 8258
rect 0 8200 1766 8256
rect 1822 8200 1827 8256
rect 0 8198 1827 8200
rect 0 8168 120 8198
rect 1761 8195 1827 8198
rect 33041 8258 33107 8261
rect 34288 8258 34408 8288
rect 33041 8256 34408 8258
rect 33041 8200 33046 8256
rect 33102 8200 34408 8256
rect 33041 8198 34408 8200
rect 33041 8195 33107 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 7946 8127 8262 8128
rect 13946 8192 14262 8193
rect 13946 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14262 8192
rect 13946 8127 14262 8128
rect 19946 8192 20262 8193
rect 19946 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20262 8192
rect 19946 8127 20262 8128
rect 25946 8192 26262 8193
rect 25946 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26262 8192
rect 25946 8127 26262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 34288 8168 34408 8198
rect 31946 8127 32262 8128
rect 0 7986 120 8016
rect 2589 7986 2655 7989
rect 0 7984 2655 7986
rect 0 7928 2594 7984
rect 2650 7928 2655 7984
rect 0 7926 2655 7928
rect 0 7896 120 7926
rect 2589 7923 2655 7926
rect 32489 7986 32555 7989
rect 34288 7986 34408 8016
rect 32489 7984 34408 7986
rect 32489 7928 32494 7984
rect 32550 7928 34408 7984
rect 32489 7926 34408 7928
rect 32489 7923 32555 7926
rect 34288 7896 34408 7926
rect 18965 7850 19031 7853
rect 2868 7848 19031 7850
rect 2868 7792 18970 7848
rect 19026 7792 19031 7848
rect 2868 7790 19031 7792
rect 0 7714 120 7744
rect 2868 7714 2928 7790
rect 18965 7787 19031 7790
rect 0 7654 2928 7714
rect 33593 7714 33659 7717
rect 34288 7714 34408 7744
rect 33593 7712 34408 7714
rect 33593 7656 33598 7712
rect 33654 7656 34408 7712
rect 33593 7654 34408 7656
rect 0 7624 120 7654
rect 33593 7651 33659 7654
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 9006 7648 9322 7649
rect 9006 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9322 7648
rect 9006 7583 9322 7584
rect 15006 7648 15322 7649
rect 15006 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15322 7648
rect 15006 7583 15322 7584
rect 21006 7648 21322 7649
rect 21006 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21322 7648
rect 21006 7583 21322 7584
rect 27006 7648 27322 7649
rect 27006 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27322 7648
rect 27006 7583 27322 7584
rect 33006 7648 33322 7649
rect 33006 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33322 7648
rect 34288 7624 34408 7654
rect 33006 7583 33322 7584
rect 0 7442 120 7472
rect 15469 7442 15535 7445
rect 0 7440 15535 7442
rect 0 7384 15474 7440
rect 15530 7384 15535 7440
rect 0 7382 15535 7384
rect 0 7352 120 7382
rect 15469 7379 15535 7382
rect 32489 7442 32555 7445
rect 34288 7442 34408 7472
rect 32489 7440 34408 7442
rect 32489 7384 32494 7440
rect 32550 7384 34408 7440
rect 32489 7382 34408 7384
rect 32489 7379 32555 7382
rect 34288 7352 34408 7382
rect 16481 7306 16547 7309
rect 1718 7304 16547 7306
rect 1718 7248 16486 7304
rect 16542 7248 16547 7304
rect 1718 7246 16547 7248
rect 0 7170 120 7200
rect 1718 7170 1778 7246
rect 16481 7243 16547 7246
rect 0 7110 1778 7170
rect 32857 7170 32923 7173
rect 34288 7170 34408 7200
rect 32857 7168 34408 7170
rect 32857 7112 32862 7168
rect 32918 7112 34408 7168
rect 32857 7110 34408 7112
rect 0 7080 120 7110
rect 32857 7107 32923 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 7946 7039 8262 7040
rect 13946 7104 14262 7105
rect 13946 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14262 7104
rect 13946 7039 14262 7040
rect 19946 7104 20262 7105
rect 19946 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20262 7104
rect 19946 7039 20262 7040
rect 25946 7104 26262 7105
rect 25946 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26262 7104
rect 25946 7039 26262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 34288 7080 34408 7110
rect 31946 7039 32262 7040
rect 0 6898 120 6928
rect 15745 6898 15811 6901
rect 0 6896 15811 6898
rect 0 6840 15750 6896
rect 15806 6840 15811 6896
rect 0 6838 15811 6840
rect 0 6808 120 6838
rect 15745 6835 15811 6838
rect 32857 6898 32923 6901
rect 34288 6898 34408 6928
rect 32857 6896 34408 6898
rect 32857 6840 32862 6896
rect 32918 6840 34408 6896
rect 32857 6838 34408 6840
rect 32857 6835 32923 6838
rect 34288 6808 34408 6838
rect 0 6626 120 6656
rect 2865 6626 2931 6629
rect 0 6624 2931 6626
rect 0 6568 2870 6624
rect 2926 6568 2931 6624
rect 0 6566 2931 6568
rect 0 6536 120 6566
rect 2865 6563 2931 6566
rect 33409 6626 33475 6629
rect 34288 6626 34408 6656
rect 33409 6624 34408 6626
rect 33409 6568 33414 6624
rect 33470 6568 34408 6624
rect 33409 6566 34408 6568
rect 33409 6563 33475 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 9006 6560 9322 6561
rect 9006 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9322 6560
rect 9006 6495 9322 6496
rect 15006 6560 15322 6561
rect 15006 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15322 6560
rect 15006 6495 15322 6496
rect 21006 6560 21322 6561
rect 21006 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21322 6560
rect 21006 6495 21322 6496
rect 27006 6560 27322 6561
rect 27006 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27322 6560
rect 27006 6495 27322 6496
rect 33006 6560 33322 6561
rect 33006 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33322 6560
rect 34288 6536 34408 6566
rect 33006 6495 33322 6496
rect 0 6354 120 6384
rect 15101 6354 15167 6357
rect 0 6352 15167 6354
rect 0 6296 15106 6352
rect 15162 6296 15167 6352
rect 0 6294 15167 6296
rect 0 6264 120 6294
rect 15101 6291 15167 6294
rect 32857 6354 32923 6357
rect 34288 6354 34408 6384
rect 32857 6352 34408 6354
rect 32857 6296 32862 6352
rect 32918 6296 34408 6352
rect 32857 6294 34408 6296
rect 32857 6291 32923 6294
rect 34288 6264 34408 6294
rect 2865 6218 2931 6221
rect 16205 6218 16271 6221
rect 2865 6216 16271 6218
rect 2865 6160 2870 6216
rect 2926 6160 16210 6216
rect 16266 6160 16271 6216
rect 2865 6158 16271 6160
rect 2865 6155 2931 6158
rect 16205 6155 16271 6158
rect 0 6082 120 6112
rect 1761 6082 1827 6085
rect 0 6080 1827 6082
rect 0 6024 1766 6080
rect 1822 6024 1827 6080
rect 0 6022 1827 6024
rect 0 5992 120 6022
rect 1761 6019 1827 6022
rect 32489 6082 32555 6085
rect 34288 6082 34408 6112
rect 32489 6080 34408 6082
rect 32489 6024 32494 6080
rect 32550 6024 34408 6080
rect 32489 6022 34408 6024
rect 32489 6019 32555 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 7946 5951 8262 5952
rect 13946 6016 14262 6017
rect 13946 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14262 6016
rect 13946 5951 14262 5952
rect 19946 6016 20262 6017
rect 19946 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20262 6016
rect 19946 5951 20262 5952
rect 25946 6016 26262 6017
rect 25946 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26262 6016
rect 25946 5951 26262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 34288 5992 34408 6022
rect 31946 5951 32262 5952
rect 0 5810 120 5840
rect 22277 5810 22343 5813
rect 0 5808 22343 5810
rect 0 5752 22282 5808
rect 22338 5752 22343 5808
rect 0 5750 22343 5752
rect 0 5720 120 5750
rect 22277 5747 22343 5750
rect 24853 5810 24919 5813
rect 25078 5810 25084 5812
rect 24853 5808 25084 5810
rect 24853 5752 24858 5808
rect 24914 5752 25084 5808
rect 24853 5750 25084 5752
rect 24853 5747 24919 5750
rect 25078 5748 25084 5750
rect 25148 5748 25154 5812
rect 32857 5810 32923 5813
rect 34288 5810 34408 5840
rect 32857 5808 34408 5810
rect 32857 5752 32862 5808
rect 32918 5752 34408 5808
rect 32857 5750 34408 5752
rect 32857 5747 32923 5750
rect 34288 5720 34408 5750
rect 1761 5674 1827 5677
rect 16389 5674 16455 5677
rect 1761 5672 16455 5674
rect 1761 5616 1766 5672
rect 1822 5616 16394 5672
rect 16450 5616 16455 5672
rect 1761 5614 16455 5616
rect 1761 5611 1827 5614
rect 16389 5611 16455 5614
rect 0 5538 120 5568
rect 2773 5538 2839 5541
rect 0 5536 2839 5538
rect 0 5480 2778 5536
rect 2834 5480 2839 5536
rect 0 5478 2839 5480
rect 0 5448 120 5478
rect 2773 5475 2839 5478
rect 33409 5538 33475 5541
rect 34288 5538 34408 5568
rect 33409 5536 34408 5538
rect 33409 5480 33414 5536
rect 33470 5480 34408 5536
rect 33409 5478 34408 5480
rect 33409 5475 33475 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 9006 5472 9322 5473
rect 9006 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9322 5472
rect 9006 5407 9322 5408
rect 15006 5472 15322 5473
rect 15006 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15322 5472
rect 15006 5407 15322 5408
rect 21006 5472 21322 5473
rect 21006 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21322 5472
rect 21006 5407 21322 5408
rect 27006 5472 27322 5473
rect 27006 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27322 5472
rect 27006 5407 27322 5408
rect 33006 5472 33322 5473
rect 33006 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33322 5472
rect 34288 5448 34408 5478
rect 33006 5407 33322 5408
rect 0 5266 120 5296
rect 2681 5266 2747 5269
rect 0 5264 2747 5266
rect 0 5208 2686 5264
rect 2742 5208 2747 5264
rect 0 5206 2747 5208
rect 0 5176 120 5206
rect 2681 5203 2747 5206
rect 15929 5266 15995 5269
rect 26693 5266 26759 5269
rect 15929 5264 26759 5266
rect 15929 5208 15934 5264
rect 15990 5208 26698 5264
rect 26754 5208 26759 5264
rect 15929 5206 26759 5208
rect 15929 5203 15995 5206
rect 26693 5203 26759 5206
rect 32857 5266 32923 5269
rect 34288 5266 34408 5296
rect 32857 5264 34408 5266
rect 32857 5208 32862 5264
rect 32918 5208 34408 5264
rect 32857 5206 34408 5208
rect 32857 5203 32923 5206
rect 34288 5176 34408 5206
rect 11053 5130 11119 5133
rect 15653 5130 15719 5133
rect 11053 5128 15719 5130
rect 11053 5072 11058 5128
rect 11114 5072 15658 5128
rect 15714 5072 15719 5128
rect 11053 5070 15719 5072
rect 11053 5067 11119 5070
rect 15653 5067 15719 5070
rect 0 4994 120 5024
rect 1301 4994 1367 4997
rect 0 4992 1367 4994
rect 0 4936 1306 4992
rect 1362 4936 1367 4992
rect 0 4934 1367 4936
rect 0 4904 120 4934
rect 1301 4931 1367 4934
rect 32489 4994 32555 4997
rect 34288 4994 34408 5024
rect 32489 4992 34408 4994
rect 32489 4936 32494 4992
rect 32550 4936 34408 4992
rect 32489 4934 34408 4936
rect 32489 4931 32555 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 13946 4928 14262 4929
rect 13946 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14262 4928
rect 13946 4863 14262 4864
rect 19946 4928 20262 4929
rect 19946 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20262 4928
rect 19946 4863 20262 4864
rect 25946 4928 26262 4929
rect 25946 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26262 4928
rect 25946 4863 26262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 34288 4904 34408 4934
rect 31946 4863 32262 4864
rect 0 4722 120 4752
rect 841 4722 907 4725
rect 0 4720 907 4722
rect 0 4664 846 4720
rect 902 4664 907 4720
rect 0 4662 907 4664
rect 0 4632 120 4662
rect 841 4659 907 4662
rect 11605 4722 11671 4725
rect 20805 4722 20871 4725
rect 11605 4720 20871 4722
rect 11605 4664 11610 4720
rect 11666 4664 20810 4720
rect 20866 4664 20871 4720
rect 11605 4662 20871 4664
rect 11605 4659 11671 4662
rect 20805 4659 20871 4662
rect 26734 4660 26740 4724
rect 26804 4722 26810 4724
rect 28441 4722 28507 4725
rect 26804 4720 28507 4722
rect 26804 4664 28446 4720
rect 28502 4664 28507 4720
rect 26804 4662 28507 4664
rect 26804 4660 26810 4662
rect 28441 4659 28507 4662
rect 32857 4722 32923 4725
rect 34288 4722 34408 4752
rect 32857 4720 34408 4722
rect 32857 4664 32862 4720
rect 32918 4664 34408 4720
rect 32857 4662 34408 4664
rect 32857 4659 32923 4662
rect 34288 4632 34408 4662
rect 1301 4586 1367 4589
rect 17125 4586 17191 4589
rect 28257 4588 28323 4589
rect 1301 4584 17191 4586
rect 1301 4528 1306 4584
rect 1362 4528 17130 4584
rect 17186 4528 17191 4584
rect 1301 4526 17191 4528
rect 1301 4523 1367 4526
rect 17125 4523 17191 4526
rect 28206 4524 28212 4588
rect 28276 4586 28323 4588
rect 28276 4584 28368 4586
rect 28318 4528 28368 4584
rect 28276 4526 28368 4528
rect 28276 4524 28323 4526
rect 28257 4523 28323 4524
rect 0 4450 120 4480
rect 1209 4450 1275 4453
rect 0 4448 1275 4450
rect 0 4392 1214 4448
rect 1270 4392 1275 4448
rect 0 4390 1275 4392
rect 0 4360 120 4390
rect 1209 4387 1275 4390
rect 33409 4450 33475 4453
rect 34288 4450 34408 4480
rect 33409 4448 34408 4450
rect 33409 4392 33414 4448
rect 33470 4392 34408 4448
rect 33409 4390 34408 4392
rect 33409 4387 33475 4390
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 9006 4384 9322 4385
rect 9006 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9322 4384
rect 9006 4319 9322 4320
rect 15006 4384 15322 4385
rect 15006 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15322 4384
rect 15006 4319 15322 4320
rect 21006 4384 21322 4385
rect 21006 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21322 4384
rect 21006 4319 21322 4320
rect 27006 4384 27322 4385
rect 27006 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27322 4384
rect 27006 4319 27322 4320
rect 33006 4384 33322 4385
rect 33006 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33322 4384
rect 34288 4360 34408 4390
rect 33006 4319 33322 4320
rect 0 4178 120 4208
rect 1117 4178 1183 4181
rect 27521 4178 27587 4181
rect 0 4176 1183 4178
rect 0 4120 1122 4176
rect 1178 4120 1183 4176
rect 0 4118 1183 4120
rect 0 4088 120 4118
rect 1117 4115 1183 4118
rect 15702 4176 27587 4178
rect 15702 4120 27526 4176
rect 27582 4120 27587 4176
rect 15702 4118 27587 4120
rect 14733 4042 14799 4045
rect 15702 4042 15762 4118
rect 27521 4115 27587 4118
rect 27654 4116 27660 4180
rect 27724 4178 27730 4180
rect 27889 4178 27955 4181
rect 27724 4176 27955 4178
rect 27724 4120 27894 4176
rect 27950 4120 27955 4176
rect 27724 4118 27955 4120
rect 27724 4116 27730 4118
rect 27889 4115 27955 4118
rect 32857 4178 32923 4181
rect 34288 4178 34408 4208
rect 32857 4176 34408 4178
rect 32857 4120 32862 4176
rect 32918 4120 34408 4176
rect 32857 4118 34408 4120
rect 32857 4115 32923 4118
rect 34288 4088 34408 4118
rect 28441 4042 28507 4045
rect 14733 4040 15762 4042
rect 14733 3984 14738 4040
rect 14794 3984 15762 4040
rect 14733 3982 15762 3984
rect 15886 4040 28507 4042
rect 15886 3984 28446 4040
rect 28502 3984 28507 4040
rect 15886 3982 28507 3984
rect 14733 3979 14799 3982
rect 0 3906 120 3936
rect 1669 3906 1735 3909
rect 0 3904 1735 3906
rect 0 3848 1674 3904
rect 1730 3848 1735 3904
rect 0 3846 1735 3848
rect 0 3816 120 3846
rect 1669 3843 1735 3846
rect 14457 3906 14523 3909
rect 15886 3906 15946 3982
rect 28441 3979 28507 3982
rect 14457 3904 15946 3906
rect 14457 3848 14462 3904
rect 14518 3848 15946 3904
rect 14457 3846 15946 3848
rect 32489 3906 32555 3909
rect 34288 3906 34408 3936
rect 32489 3904 34408 3906
rect 32489 3848 32494 3904
rect 32550 3848 34408 3904
rect 32489 3846 34408 3848
rect 14457 3843 14523 3846
rect 32489 3843 32555 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 13946 3840 14262 3841
rect 13946 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14262 3840
rect 13946 3775 14262 3776
rect 19946 3840 20262 3841
rect 19946 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20262 3840
rect 19946 3775 20262 3776
rect 25946 3840 26262 3841
rect 25946 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26262 3840
rect 25946 3775 26262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 34288 3816 34408 3846
rect 31946 3775 32262 3776
rect 26325 3770 26391 3773
rect 31661 3770 31727 3773
rect 26325 3768 31727 3770
rect 26325 3712 26330 3768
rect 26386 3712 31666 3768
rect 31722 3712 31727 3768
rect 26325 3710 31727 3712
rect 26325 3707 26391 3710
rect 31661 3707 31727 3710
rect 0 3634 120 3664
rect 20713 3634 20779 3637
rect 0 3632 20779 3634
rect 0 3576 20718 3632
rect 20774 3576 20779 3632
rect 0 3574 20779 3576
rect 0 3544 120 3574
rect 20713 3571 20779 3574
rect 24761 3634 24827 3637
rect 30373 3634 30439 3637
rect 24761 3632 30439 3634
rect 24761 3576 24766 3632
rect 24822 3576 30378 3632
rect 30434 3576 30439 3632
rect 24761 3574 30439 3576
rect 24761 3571 24827 3574
rect 30373 3571 30439 3574
rect 32857 3634 32923 3637
rect 34288 3634 34408 3664
rect 32857 3632 34408 3634
rect 32857 3576 32862 3632
rect 32918 3576 34408 3632
rect 32857 3574 34408 3576
rect 32857 3571 32923 3574
rect 34288 3544 34408 3574
rect 2497 3498 2563 3501
rect 16757 3498 16823 3501
rect 2497 3496 16823 3498
rect 2497 3440 2502 3496
rect 2558 3440 16762 3496
rect 16818 3440 16823 3496
rect 2497 3438 16823 3440
rect 2497 3435 2563 3438
rect 16757 3435 16823 3438
rect 24117 3498 24183 3501
rect 28257 3498 28323 3501
rect 24117 3496 28323 3498
rect 24117 3440 24122 3496
rect 24178 3440 28262 3496
rect 28318 3440 28323 3496
rect 24117 3438 28323 3440
rect 24117 3435 24183 3438
rect 28257 3435 28323 3438
rect 0 3362 120 3392
rect 2865 3362 2931 3365
rect 0 3360 2931 3362
rect 0 3304 2870 3360
rect 2926 3304 2931 3360
rect 0 3302 2931 3304
rect 0 3272 120 3302
rect 2865 3299 2931 3302
rect 21633 3362 21699 3365
rect 22185 3362 22251 3365
rect 21633 3360 22251 3362
rect 21633 3304 21638 3360
rect 21694 3304 22190 3360
rect 22246 3304 22251 3360
rect 21633 3302 22251 3304
rect 21633 3299 21699 3302
rect 22185 3299 22251 3302
rect 33409 3362 33475 3365
rect 34288 3362 34408 3392
rect 33409 3360 34408 3362
rect 33409 3304 33414 3360
rect 33470 3304 34408 3360
rect 33409 3302 34408 3304
rect 33409 3299 33475 3302
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 9006 3296 9322 3297
rect 9006 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9322 3296
rect 9006 3231 9322 3232
rect 15006 3296 15322 3297
rect 15006 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15322 3296
rect 15006 3231 15322 3232
rect 21006 3296 21322 3297
rect 21006 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21322 3296
rect 21006 3231 21322 3232
rect 27006 3296 27322 3297
rect 27006 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27322 3296
rect 27006 3231 27322 3232
rect 33006 3296 33322 3297
rect 33006 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33322 3296
rect 34288 3272 34408 3302
rect 33006 3231 33322 3232
rect 0 3090 120 3120
rect 23565 3090 23631 3093
rect 0 3088 23631 3090
rect 0 3032 23570 3088
rect 23626 3032 23631 3088
rect 0 3030 23631 3032
rect 0 3000 120 3030
rect 23565 3027 23631 3030
rect 24577 3090 24643 3093
rect 28441 3090 28507 3093
rect 24577 3088 28507 3090
rect 24577 3032 24582 3088
rect 24638 3032 28446 3088
rect 28502 3032 28507 3088
rect 24577 3030 28507 3032
rect 24577 3027 24643 3030
rect 28441 3027 28507 3030
rect 32857 3090 32923 3093
rect 34288 3090 34408 3120
rect 32857 3088 34408 3090
rect 32857 3032 32862 3088
rect 32918 3032 34408 3088
rect 32857 3030 34408 3032
rect 32857 3027 32923 3030
rect 34288 3000 34408 3030
rect 2865 2954 2931 2957
rect 24853 2954 24919 2957
rect 2865 2952 24919 2954
rect 2865 2896 2870 2952
rect 2926 2896 24858 2952
rect 24914 2896 24919 2952
rect 2865 2894 24919 2896
rect 2865 2891 2931 2894
rect 24853 2891 24919 2894
rect 25630 2892 25636 2956
rect 25700 2954 25706 2956
rect 27797 2954 27863 2957
rect 25700 2952 27863 2954
rect 25700 2896 27802 2952
rect 27858 2896 27863 2952
rect 25700 2894 27863 2896
rect 25700 2892 25706 2894
rect 27797 2891 27863 2894
rect 0 2818 120 2848
rect 1301 2818 1367 2821
rect 0 2816 1367 2818
rect 0 2760 1306 2816
rect 1362 2760 1367 2816
rect 0 2758 1367 2760
rect 0 2728 120 2758
rect 1301 2755 1367 2758
rect 14825 2818 14891 2821
rect 16021 2818 16087 2821
rect 14825 2816 16087 2818
rect 14825 2760 14830 2816
rect 14886 2760 16026 2816
rect 16082 2760 16087 2816
rect 14825 2758 16087 2760
rect 14825 2755 14891 2758
rect 16021 2755 16087 2758
rect 32489 2818 32555 2821
rect 34288 2818 34408 2848
rect 32489 2816 34408 2818
rect 32489 2760 32494 2816
rect 32550 2760 34408 2816
rect 32489 2758 34408 2760
rect 32489 2755 32555 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 13946 2752 14262 2753
rect 13946 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14262 2752
rect 13946 2687 14262 2688
rect 19946 2752 20262 2753
rect 19946 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20262 2752
rect 19946 2687 20262 2688
rect 25946 2752 26262 2753
rect 25946 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26262 2752
rect 25946 2687 26262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 34288 2728 34408 2758
rect 31946 2687 32262 2688
rect 23013 2682 23079 2685
rect 25497 2682 25563 2685
rect 23013 2680 25563 2682
rect 23013 2624 23018 2680
rect 23074 2624 25502 2680
rect 25558 2624 25563 2680
rect 23013 2622 25563 2624
rect 23013 2619 23079 2622
rect 25497 2619 25563 2622
rect 0 2546 120 2576
rect 23381 2546 23447 2549
rect 0 2544 23447 2546
rect 0 2488 23386 2544
rect 23442 2488 23447 2544
rect 0 2486 23447 2488
rect 0 2456 120 2486
rect 23381 2483 23447 2486
rect 23933 2546 23999 2549
rect 25773 2546 25839 2549
rect 23933 2544 25839 2546
rect 23933 2488 23938 2544
rect 23994 2488 25778 2544
rect 25834 2488 25839 2544
rect 23933 2486 25839 2488
rect 23933 2483 23999 2486
rect 25773 2483 25839 2486
rect 26049 2546 26115 2549
rect 26734 2546 26740 2548
rect 26049 2544 26740 2546
rect 26049 2488 26054 2544
rect 26110 2488 26740 2544
rect 26049 2486 26740 2488
rect 26049 2483 26115 2486
rect 26734 2484 26740 2486
rect 26804 2484 26810 2548
rect 32857 2546 32923 2549
rect 34288 2546 34408 2576
rect 32857 2544 34408 2546
rect 32857 2488 32862 2544
rect 32918 2488 34408 2544
rect 32857 2486 34408 2488
rect 32857 2483 32923 2486
rect 34288 2456 34408 2486
rect 12433 2410 12499 2413
rect 26877 2410 26943 2413
rect 12433 2408 26943 2410
rect 12433 2352 12438 2408
rect 12494 2352 26882 2408
rect 26938 2352 26943 2408
rect 12433 2350 26943 2352
rect 12433 2347 12499 2350
rect 26877 2347 26943 2350
rect 0 2274 120 2304
rect 2865 2274 2931 2277
rect 0 2272 2931 2274
rect 0 2216 2870 2272
rect 2926 2216 2931 2272
rect 0 2214 2931 2216
rect 0 2184 120 2214
rect 2865 2211 2931 2214
rect 33409 2274 33475 2277
rect 34288 2274 34408 2304
rect 33409 2272 34408 2274
rect 33409 2216 33414 2272
rect 33470 2216 34408 2272
rect 33409 2214 34408 2216
rect 33409 2211 33475 2214
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 9006 2208 9322 2209
rect 9006 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9322 2208
rect 9006 2143 9322 2144
rect 15006 2208 15322 2209
rect 15006 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15322 2208
rect 15006 2143 15322 2144
rect 21006 2208 21322 2209
rect 21006 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21322 2208
rect 21006 2143 21322 2144
rect 27006 2208 27322 2209
rect 27006 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27322 2208
rect 27006 2143 27322 2144
rect 33006 2208 33322 2209
rect 33006 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33322 2208
rect 34288 2184 34408 2214
rect 33006 2143 33322 2144
rect 9857 2138 9923 2141
rect 13813 2138 13879 2141
rect 9857 2136 13879 2138
rect 9857 2080 9862 2136
rect 9918 2080 13818 2136
rect 13874 2080 13879 2136
rect 9857 2078 13879 2080
rect 9857 2075 9923 2078
rect 13813 2075 13879 2078
rect 0 2002 120 2032
rect 21909 2002 21975 2005
rect 0 2000 21975 2002
rect 0 1944 21914 2000
rect 21970 1944 21975 2000
rect 0 1942 21975 1944
rect 0 1912 120 1942
rect 21909 1939 21975 1942
rect 31109 2002 31175 2005
rect 34288 2002 34408 2032
rect 31109 2000 34408 2002
rect 31109 1944 31114 2000
rect 31170 1944 34408 2000
rect 31109 1942 34408 1944
rect 31109 1939 31175 1942
rect 34288 1912 34408 1942
rect 2865 1866 2931 1869
rect 17493 1866 17559 1869
rect 2865 1864 17559 1866
rect 2865 1808 2870 1864
rect 2926 1808 17498 1864
rect 17554 1808 17559 1864
rect 2865 1806 17559 1808
rect 2865 1803 2931 1806
rect 17493 1803 17559 1806
rect 19701 1866 19767 1869
rect 25313 1866 25379 1869
rect 19701 1864 25379 1866
rect 19701 1808 19706 1864
rect 19762 1808 25318 1864
rect 25374 1808 25379 1864
rect 19701 1806 25379 1808
rect 19701 1803 19767 1806
rect 25313 1803 25379 1806
rect 0 1730 120 1760
rect 16757 1730 16823 1733
rect 0 1728 16823 1730
rect 0 1672 16762 1728
rect 16818 1672 16823 1728
rect 0 1670 16823 1672
rect 0 1640 120 1670
rect 16757 1667 16823 1670
rect 32397 1730 32463 1733
rect 34288 1730 34408 1760
rect 32397 1728 34408 1730
rect 32397 1672 32402 1728
rect 32458 1672 34408 1728
rect 32397 1670 34408 1672
rect 32397 1667 32463 1670
rect 34288 1640 34408 1670
rect 0 1458 120 1488
rect 19425 1458 19491 1461
rect 0 1456 19491 1458
rect 0 1400 19430 1456
rect 19486 1400 19491 1456
rect 0 1398 19491 1400
rect 0 1368 120 1398
rect 19425 1395 19491 1398
rect 27521 1458 27587 1461
rect 30465 1458 30531 1461
rect 27521 1456 30531 1458
rect 27521 1400 27526 1456
rect 27582 1400 30470 1456
rect 30526 1400 30531 1456
rect 27521 1398 30531 1400
rect 27521 1395 27587 1398
rect 30465 1395 30531 1398
rect 31477 1458 31543 1461
rect 34288 1458 34408 1488
rect 31477 1456 34408 1458
rect 31477 1400 31482 1456
rect 31538 1400 34408 1456
rect 31477 1398 34408 1400
rect 31477 1395 31543 1398
rect 34288 1368 34408 1398
rect 4521 1322 4587 1325
rect 7465 1322 7531 1325
rect 4521 1320 7531 1322
rect 4521 1264 4526 1320
rect 4582 1264 7470 1320
rect 7526 1264 7531 1320
rect 4521 1262 7531 1264
rect 4521 1259 4587 1262
rect 7465 1259 7531 1262
rect 25589 1322 25655 1325
rect 26969 1322 27035 1325
rect 25589 1320 27035 1322
rect 25589 1264 25594 1320
rect 25650 1264 26974 1320
rect 27030 1264 27035 1320
rect 25589 1262 27035 1264
rect 25589 1259 25655 1262
rect 26969 1259 27035 1262
rect 0 1186 120 1216
rect 17677 1186 17743 1189
rect 0 1184 17743 1186
rect 0 1128 17682 1184
rect 17738 1128 17743 1184
rect 0 1126 17743 1128
rect 0 1096 120 1126
rect 17677 1123 17743 1126
rect 31845 1186 31911 1189
rect 34288 1186 34408 1216
rect 31845 1184 34408 1186
rect 31845 1128 31850 1184
rect 31906 1128 34408 1184
rect 31845 1126 34408 1128
rect 31845 1123 31911 1126
rect 34288 1096 34408 1126
rect 13721 642 13787 645
rect 25630 642 25636 644
rect 13721 640 25636 642
rect 13721 584 13726 640
rect 13782 584 25636 640
rect 13721 582 25636 584
rect 13721 579 13787 582
rect 25630 580 25636 582
rect 25700 580 25706 644
rect 13537 506 13603 509
rect 28206 506 28212 508
rect 13537 504 28212 506
rect 13537 448 13542 504
rect 13598 448 28212 504
rect 13537 446 28212 448
rect 13537 443 13603 446
rect 28206 444 28212 446
rect 28276 444 28282 508
rect 13353 370 13419 373
rect 26877 370 26943 373
rect 13353 368 26943 370
rect 13353 312 13358 368
rect 13414 312 26882 368
rect 26938 312 26943 368
rect 13353 310 26943 312
rect 13353 307 13419 310
rect 26877 307 26943 310
rect 13905 234 13971 237
rect 27654 234 27660 236
rect 13905 232 27660 234
rect 13905 176 13910 232
rect 13966 176 27660 232
rect 13905 174 27660 176
rect 13905 171 13971 174
rect 27654 172 27660 174
rect 27724 172 27730 236
rect 4889 98 4955 101
rect 7649 98 7715 101
rect 25129 100 25195 101
rect 4889 96 7715 98
rect 4889 40 4894 96
rect 4950 40 7654 96
rect 7710 40 7715 96
rect 4889 38 7715 40
rect 4889 35 4955 38
rect 7649 35 7715 38
rect 25078 36 25084 100
rect 25148 98 25195 100
rect 25405 98 25471 101
rect 26601 98 26667 101
rect 25148 96 25240 98
rect 25190 40 25240 96
rect 25148 38 25240 40
rect 25405 96 26667 98
rect 25405 40 25410 96
rect 25466 40 26606 96
rect 26662 40 26667 96
rect 25405 38 26667 40
rect 25148 36 25195 38
rect 25129 35 25195 36
rect 25405 35 25471 38
rect 26601 35 26667 38
<< via3 >>
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 9172 8732 9236 8736
rect 9172 8676 9176 8732
rect 9176 8676 9232 8732
rect 9232 8676 9236 8732
rect 9172 8672 9236 8676
rect 9252 8732 9316 8736
rect 9252 8676 9256 8732
rect 9256 8676 9312 8732
rect 9312 8676 9316 8732
rect 9252 8672 9316 8676
rect 15012 8732 15076 8736
rect 15012 8676 15016 8732
rect 15016 8676 15072 8732
rect 15072 8676 15076 8732
rect 15012 8672 15076 8676
rect 15092 8732 15156 8736
rect 15092 8676 15096 8732
rect 15096 8676 15152 8732
rect 15152 8676 15156 8732
rect 15092 8672 15156 8676
rect 15172 8732 15236 8736
rect 15172 8676 15176 8732
rect 15176 8676 15232 8732
rect 15232 8676 15236 8732
rect 15172 8672 15236 8676
rect 15252 8732 15316 8736
rect 15252 8676 15256 8732
rect 15256 8676 15312 8732
rect 15312 8676 15316 8732
rect 15252 8672 15316 8676
rect 21012 8732 21076 8736
rect 21012 8676 21016 8732
rect 21016 8676 21072 8732
rect 21072 8676 21076 8732
rect 21012 8672 21076 8676
rect 21092 8732 21156 8736
rect 21092 8676 21096 8732
rect 21096 8676 21152 8732
rect 21152 8676 21156 8732
rect 21092 8672 21156 8676
rect 21172 8732 21236 8736
rect 21172 8676 21176 8732
rect 21176 8676 21232 8732
rect 21232 8676 21236 8732
rect 21172 8672 21236 8676
rect 21252 8732 21316 8736
rect 21252 8676 21256 8732
rect 21256 8676 21312 8732
rect 21312 8676 21316 8732
rect 21252 8672 21316 8676
rect 27012 8732 27076 8736
rect 27012 8676 27016 8732
rect 27016 8676 27072 8732
rect 27072 8676 27076 8732
rect 27012 8672 27076 8676
rect 27092 8732 27156 8736
rect 27092 8676 27096 8732
rect 27096 8676 27152 8732
rect 27152 8676 27156 8732
rect 27092 8672 27156 8676
rect 27172 8732 27236 8736
rect 27172 8676 27176 8732
rect 27176 8676 27232 8732
rect 27232 8676 27236 8732
rect 27172 8672 27236 8676
rect 27252 8732 27316 8736
rect 27252 8676 27256 8732
rect 27256 8676 27312 8732
rect 27312 8676 27316 8732
rect 27252 8672 27316 8676
rect 33012 8732 33076 8736
rect 33012 8676 33016 8732
rect 33016 8676 33072 8732
rect 33072 8676 33076 8732
rect 33012 8672 33076 8676
rect 33092 8732 33156 8736
rect 33092 8676 33096 8732
rect 33096 8676 33152 8732
rect 33152 8676 33156 8732
rect 33092 8672 33156 8676
rect 33172 8732 33236 8736
rect 33172 8676 33176 8732
rect 33176 8676 33232 8732
rect 33232 8676 33236 8732
rect 33172 8672 33236 8676
rect 33252 8732 33316 8736
rect 33252 8676 33256 8732
rect 33256 8676 33312 8732
rect 33312 8676 33316 8732
rect 33252 8672 33316 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 13952 8188 14016 8192
rect 13952 8132 13956 8188
rect 13956 8132 14012 8188
rect 14012 8132 14016 8188
rect 13952 8128 14016 8132
rect 14032 8188 14096 8192
rect 14032 8132 14036 8188
rect 14036 8132 14092 8188
rect 14092 8132 14096 8188
rect 14032 8128 14096 8132
rect 14112 8188 14176 8192
rect 14112 8132 14116 8188
rect 14116 8132 14172 8188
rect 14172 8132 14176 8188
rect 14112 8128 14176 8132
rect 14192 8188 14256 8192
rect 14192 8132 14196 8188
rect 14196 8132 14252 8188
rect 14252 8132 14256 8188
rect 14192 8128 14256 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 20192 8188 20256 8192
rect 20192 8132 20196 8188
rect 20196 8132 20252 8188
rect 20252 8132 20256 8188
rect 20192 8128 20256 8132
rect 25952 8188 26016 8192
rect 25952 8132 25956 8188
rect 25956 8132 26012 8188
rect 26012 8132 26016 8188
rect 25952 8128 26016 8132
rect 26032 8188 26096 8192
rect 26032 8132 26036 8188
rect 26036 8132 26092 8188
rect 26092 8132 26096 8188
rect 26032 8128 26096 8132
rect 26112 8188 26176 8192
rect 26112 8132 26116 8188
rect 26116 8132 26172 8188
rect 26172 8132 26176 8188
rect 26112 8128 26176 8132
rect 26192 8188 26256 8192
rect 26192 8132 26196 8188
rect 26196 8132 26252 8188
rect 26252 8132 26256 8188
rect 26192 8128 26256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 9172 7644 9236 7648
rect 9172 7588 9176 7644
rect 9176 7588 9232 7644
rect 9232 7588 9236 7644
rect 9172 7584 9236 7588
rect 9252 7644 9316 7648
rect 9252 7588 9256 7644
rect 9256 7588 9312 7644
rect 9312 7588 9316 7644
rect 9252 7584 9316 7588
rect 15012 7644 15076 7648
rect 15012 7588 15016 7644
rect 15016 7588 15072 7644
rect 15072 7588 15076 7644
rect 15012 7584 15076 7588
rect 15092 7644 15156 7648
rect 15092 7588 15096 7644
rect 15096 7588 15152 7644
rect 15152 7588 15156 7644
rect 15092 7584 15156 7588
rect 15172 7644 15236 7648
rect 15172 7588 15176 7644
rect 15176 7588 15232 7644
rect 15232 7588 15236 7644
rect 15172 7584 15236 7588
rect 15252 7644 15316 7648
rect 15252 7588 15256 7644
rect 15256 7588 15312 7644
rect 15312 7588 15316 7644
rect 15252 7584 15316 7588
rect 21012 7644 21076 7648
rect 21012 7588 21016 7644
rect 21016 7588 21072 7644
rect 21072 7588 21076 7644
rect 21012 7584 21076 7588
rect 21092 7644 21156 7648
rect 21092 7588 21096 7644
rect 21096 7588 21152 7644
rect 21152 7588 21156 7644
rect 21092 7584 21156 7588
rect 21172 7644 21236 7648
rect 21172 7588 21176 7644
rect 21176 7588 21232 7644
rect 21232 7588 21236 7644
rect 21172 7584 21236 7588
rect 21252 7644 21316 7648
rect 21252 7588 21256 7644
rect 21256 7588 21312 7644
rect 21312 7588 21316 7644
rect 21252 7584 21316 7588
rect 27012 7644 27076 7648
rect 27012 7588 27016 7644
rect 27016 7588 27072 7644
rect 27072 7588 27076 7644
rect 27012 7584 27076 7588
rect 27092 7644 27156 7648
rect 27092 7588 27096 7644
rect 27096 7588 27152 7644
rect 27152 7588 27156 7644
rect 27092 7584 27156 7588
rect 27172 7644 27236 7648
rect 27172 7588 27176 7644
rect 27176 7588 27232 7644
rect 27232 7588 27236 7644
rect 27172 7584 27236 7588
rect 27252 7644 27316 7648
rect 27252 7588 27256 7644
rect 27256 7588 27312 7644
rect 27312 7588 27316 7644
rect 27252 7584 27316 7588
rect 33012 7644 33076 7648
rect 33012 7588 33016 7644
rect 33016 7588 33072 7644
rect 33072 7588 33076 7644
rect 33012 7584 33076 7588
rect 33092 7644 33156 7648
rect 33092 7588 33096 7644
rect 33096 7588 33152 7644
rect 33152 7588 33156 7644
rect 33092 7584 33156 7588
rect 33172 7644 33236 7648
rect 33172 7588 33176 7644
rect 33176 7588 33232 7644
rect 33232 7588 33236 7644
rect 33172 7584 33236 7588
rect 33252 7644 33316 7648
rect 33252 7588 33256 7644
rect 33256 7588 33312 7644
rect 33312 7588 33316 7644
rect 33252 7584 33316 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 13952 7100 14016 7104
rect 13952 7044 13956 7100
rect 13956 7044 14012 7100
rect 14012 7044 14016 7100
rect 13952 7040 14016 7044
rect 14032 7100 14096 7104
rect 14032 7044 14036 7100
rect 14036 7044 14092 7100
rect 14092 7044 14096 7100
rect 14032 7040 14096 7044
rect 14112 7100 14176 7104
rect 14112 7044 14116 7100
rect 14116 7044 14172 7100
rect 14172 7044 14176 7100
rect 14112 7040 14176 7044
rect 14192 7100 14256 7104
rect 14192 7044 14196 7100
rect 14196 7044 14252 7100
rect 14252 7044 14256 7100
rect 14192 7040 14256 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 20192 7100 20256 7104
rect 20192 7044 20196 7100
rect 20196 7044 20252 7100
rect 20252 7044 20256 7100
rect 20192 7040 20256 7044
rect 25952 7100 26016 7104
rect 25952 7044 25956 7100
rect 25956 7044 26012 7100
rect 26012 7044 26016 7100
rect 25952 7040 26016 7044
rect 26032 7100 26096 7104
rect 26032 7044 26036 7100
rect 26036 7044 26092 7100
rect 26092 7044 26096 7100
rect 26032 7040 26096 7044
rect 26112 7100 26176 7104
rect 26112 7044 26116 7100
rect 26116 7044 26172 7100
rect 26172 7044 26176 7100
rect 26112 7040 26176 7044
rect 26192 7100 26256 7104
rect 26192 7044 26196 7100
rect 26196 7044 26252 7100
rect 26252 7044 26256 7100
rect 26192 7040 26256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 9172 6556 9236 6560
rect 9172 6500 9176 6556
rect 9176 6500 9232 6556
rect 9232 6500 9236 6556
rect 9172 6496 9236 6500
rect 9252 6556 9316 6560
rect 9252 6500 9256 6556
rect 9256 6500 9312 6556
rect 9312 6500 9316 6556
rect 9252 6496 9316 6500
rect 15012 6556 15076 6560
rect 15012 6500 15016 6556
rect 15016 6500 15072 6556
rect 15072 6500 15076 6556
rect 15012 6496 15076 6500
rect 15092 6556 15156 6560
rect 15092 6500 15096 6556
rect 15096 6500 15152 6556
rect 15152 6500 15156 6556
rect 15092 6496 15156 6500
rect 15172 6556 15236 6560
rect 15172 6500 15176 6556
rect 15176 6500 15232 6556
rect 15232 6500 15236 6556
rect 15172 6496 15236 6500
rect 15252 6556 15316 6560
rect 15252 6500 15256 6556
rect 15256 6500 15312 6556
rect 15312 6500 15316 6556
rect 15252 6496 15316 6500
rect 21012 6556 21076 6560
rect 21012 6500 21016 6556
rect 21016 6500 21072 6556
rect 21072 6500 21076 6556
rect 21012 6496 21076 6500
rect 21092 6556 21156 6560
rect 21092 6500 21096 6556
rect 21096 6500 21152 6556
rect 21152 6500 21156 6556
rect 21092 6496 21156 6500
rect 21172 6556 21236 6560
rect 21172 6500 21176 6556
rect 21176 6500 21232 6556
rect 21232 6500 21236 6556
rect 21172 6496 21236 6500
rect 21252 6556 21316 6560
rect 21252 6500 21256 6556
rect 21256 6500 21312 6556
rect 21312 6500 21316 6556
rect 21252 6496 21316 6500
rect 27012 6556 27076 6560
rect 27012 6500 27016 6556
rect 27016 6500 27072 6556
rect 27072 6500 27076 6556
rect 27012 6496 27076 6500
rect 27092 6556 27156 6560
rect 27092 6500 27096 6556
rect 27096 6500 27152 6556
rect 27152 6500 27156 6556
rect 27092 6496 27156 6500
rect 27172 6556 27236 6560
rect 27172 6500 27176 6556
rect 27176 6500 27232 6556
rect 27232 6500 27236 6556
rect 27172 6496 27236 6500
rect 27252 6556 27316 6560
rect 27252 6500 27256 6556
rect 27256 6500 27312 6556
rect 27312 6500 27316 6556
rect 27252 6496 27316 6500
rect 33012 6556 33076 6560
rect 33012 6500 33016 6556
rect 33016 6500 33072 6556
rect 33072 6500 33076 6556
rect 33012 6496 33076 6500
rect 33092 6556 33156 6560
rect 33092 6500 33096 6556
rect 33096 6500 33152 6556
rect 33152 6500 33156 6556
rect 33092 6496 33156 6500
rect 33172 6556 33236 6560
rect 33172 6500 33176 6556
rect 33176 6500 33232 6556
rect 33232 6500 33236 6556
rect 33172 6496 33236 6500
rect 33252 6556 33316 6560
rect 33252 6500 33256 6556
rect 33256 6500 33312 6556
rect 33312 6500 33316 6556
rect 33252 6496 33316 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 13952 6012 14016 6016
rect 13952 5956 13956 6012
rect 13956 5956 14012 6012
rect 14012 5956 14016 6012
rect 13952 5952 14016 5956
rect 14032 6012 14096 6016
rect 14032 5956 14036 6012
rect 14036 5956 14092 6012
rect 14092 5956 14096 6012
rect 14032 5952 14096 5956
rect 14112 6012 14176 6016
rect 14112 5956 14116 6012
rect 14116 5956 14172 6012
rect 14172 5956 14176 6012
rect 14112 5952 14176 5956
rect 14192 6012 14256 6016
rect 14192 5956 14196 6012
rect 14196 5956 14252 6012
rect 14252 5956 14256 6012
rect 14192 5952 14256 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 20192 6012 20256 6016
rect 20192 5956 20196 6012
rect 20196 5956 20252 6012
rect 20252 5956 20256 6012
rect 20192 5952 20256 5956
rect 25952 6012 26016 6016
rect 25952 5956 25956 6012
rect 25956 5956 26012 6012
rect 26012 5956 26016 6012
rect 25952 5952 26016 5956
rect 26032 6012 26096 6016
rect 26032 5956 26036 6012
rect 26036 5956 26092 6012
rect 26092 5956 26096 6012
rect 26032 5952 26096 5956
rect 26112 6012 26176 6016
rect 26112 5956 26116 6012
rect 26116 5956 26172 6012
rect 26172 5956 26176 6012
rect 26112 5952 26176 5956
rect 26192 6012 26256 6016
rect 26192 5956 26196 6012
rect 26196 5956 26252 6012
rect 26252 5956 26256 6012
rect 26192 5952 26256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 25084 5748 25148 5812
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 9172 5468 9236 5472
rect 9172 5412 9176 5468
rect 9176 5412 9232 5468
rect 9232 5412 9236 5468
rect 9172 5408 9236 5412
rect 9252 5468 9316 5472
rect 9252 5412 9256 5468
rect 9256 5412 9312 5468
rect 9312 5412 9316 5468
rect 9252 5408 9316 5412
rect 15012 5468 15076 5472
rect 15012 5412 15016 5468
rect 15016 5412 15072 5468
rect 15072 5412 15076 5468
rect 15012 5408 15076 5412
rect 15092 5468 15156 5472
rect 15092 5412 15096 5468
rect 15096 5412 15152 5468
rect 15152 5412 15156 5468
rect 15092 5408 15156 5412
rect 15172 5468 15236 5472
rect 15172 5412 15176 5468
rect 15176 5412 15232 5468
rect 15232 5412 15236 5468
rect 15172 5408 15236 5412
rect 15252 5468 15316 5472
rect 15252 5412 15256 5468
rect 15256 5412 15312 5468
rect 15312 5412 15316 5468
rect 15252 5408 15316 5412
rect 21012 5468 21076 5472
rect 21012 5412 21016 5468
rect 21016 5412 21072 5468
rect 21072 5412 21076 5468
rect 21012 5408 21076 5412
rect 21092 5468 21156 5472
rect 21092 5412 21096 5468
rect 21096 5412 21152 5468
rect 21152 5412 21156 5468
rect 21092 5408 21156 5412
rect 21172 5468 21236 5472
rect 21172 5412 21176 5468
rect 21176 5412 21232 5468
rect 21232 5412 21236 5468
rect 21172 5408 21236 5412
rect 21252 5468 21316 5472
rect 21252 5412 21256 5468
rect 21256 5412 21312 5468
rect 21312 5412 21316 5468
rect 21252 5408 21316 5412
rect 27012 5468 27076 5472
rect 27012 5412 27016 5468
rect 27016 5412 27072 5468
rect 27072 5412 27076 5468
rect 27012 5408 27076 5412
rect 27092 5468 27156 5472
rect 27092 5412 27096 5468
rect 27096 5412 27152 5468
rect 27152 5412 27156 5468
rect 27092 5408 27156 5412
rect 27172 5468 27236 5472
rect 27172 5412 27176 5468
rect 27176 5412 27232 5468
rect 27232 5412 27236 5468
rect 27172 5408 27236 5412
rect 27252 5468 27316 5472
rect 27252 5412 27256 5468
rect 27256 5412 27312 5468
rect 27312 5412 27316 5468
rect 27252 5408 27316 5412
rect 33012 5468 33076 5472
rect 33012 5412 33016 5468
rect 33016 5412 33072 5468
rect 33072 5412 33076 5468
rect 33012 5408 33076 5412
rect 33092 5468 33156 5472
rect 33092 5412 33096 5468
rect 33096 5412 33152 5468
rect 33152 5412 33156 5468
rect 33092 5408 33156 5412
rect 33172 5468 33236 5472
rect 33172 5412 33176 5468
rect 33176 5412 33232 5468
rect 33232 5412 33236 5468
rect 33172 5408 33236 5412
rect 33252 5468 33316 5472
rect 33252 5412 33256 5468
rect 33256 5412 33312 5468
rect 33312 5412 33316 5468
rect 33252 5408 33316 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 13952 4924 14016 4928
rect 13952 4868 13956 4924
rect 13956 4868 14012 4924
rect 14012 4868 14016 4924
rect 13952 4864 14016 4868
rect 14032 4924 14096 4928
rect 14032 4868 14036 4924
rect 14036 4868 14092 4924
rect 14092 4868 14096 4924
rect 14032 4864 14096 4868
rect 14112 4924 14176 4928
rect 14112 4868 14116 4924
rect 14116 4868 14172 4924
rect 14172 4868 14176 4924
rect 14112 4864 14176 4868
rect 14192 4924 14256 4928
rect 14192 4868 14196 4924
rect 14196 4868 14252 4924
rect 14252 4868 14256 4924
rect 14192 4864 14256 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 20192 4924 20256 4928
rect 20192 4868 20196 4924
rect 20196 4868 20252 4924
rect 20252 4868 20256 4924
rect 20192 4864 20256 4868
rect 25952 4924 26016 4928
rect 25952 4868 25956 4924
rect 25956 4868 26012 4924
rect 26012 4868 26016 4924
rect 25952 4864 26016 4868
rect 26032 4924 26096 4928
rect 26032 4868 26036 4924
rect 26036 4868 26092 4924
rect 26092 4868 26096 4924
rect 26032 4864 26096 4868
rect 26112 4924 26176 4928
rect 26112 4868 26116 4924
rect 26116 4868 26172 4924
rect 26172 4868 26176 4924
rect 26112 4864 26176 4868
rect 26192 4924 26256 4928
rect 26192 4868 26196 4924
rect 26196 4868 26252 4924
rect 26252 4868 26256 4924
rect 26192 4864 26256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 26740 4660 26804 4724
rect 28212 4584 28276 4588
rect 28212 4528 28262 4584
rect 28262 4528 28276 4584
rect 28212 4524 28276 4528
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 9172 4380 9236 4384
rect 9172 4324 9176 4380
rect 9176 4324 9232 4380
rect 9232 4324 9236 4380
rect 9172 4320 9236 4324
rect 9252 4380 9316 4384
rect 9252 4324 9256 4380
rect 9256 4324 9312 4380
rect 9312 4324 9316 4380
rect 9252 4320 9316 4324
rect 15012 4380 15076 4384
rect 15012 4324 15016 4380
rect 15016 4324 15072 4380
rect 15072 4324 15076 4380
rect 15012 4320 15076 4324
rect 15092 4380 15156 4384
rect 15092 4324 15096 4380
rect 15096 4324 15152 4380
rect 15152 4324 15156 4380
rect 15092 4320 15156 4324
rect 15172 4380 15236 4384
rect 15172 4324 15176 4380
rect 15176 4324 15232 4380
rect 15232 4324 15236 4380
rect 15172 4320 15236 4324
rect 15252 4380 15316 4384
rect 15252 4324 15256 4380
rect 15256 4324 15312 4380
rect 15312 4324 15316 4380
rect 15252 4320 15316 4324
rect 21012 4380 21076 4384
rect 21012 4324 21016 4380
rect 21016 4324 21072 4380
rect 21072 4324 21076 4380
rect 21012 4320 21076 4324
rect 21092 4380 21156 4384
rect 21092 4324 21096 4380
rect 21096 4324 21152 4380
rect 21152 4324 21156 4380
rect 21092 4320 21156 4324
rect 21172 4380 21236 4384
rect 21172 4324 21176 4380
rect 21176 4324 21232 4380
rect 21232 4324 21236 4380
rect 21172 4320 21236 4324
rect 21252 4380 21316 4384
rect 21252 4324 21256 4380
rect 21256 4324 21312 4380
rect 21312 4324 21316 4380
rect 21252 4320 21316 4324
rect 27012 4380 27076 4384
rect 27012 4324 27016 4380
rect 27016 4324 27072 4380
rect 27072 4324 27076 4380
rect 27012 4320 27076 4324
rect 27092 4380 27156 4384
rect 27092 4324 27096 4380
rect 27096 4324 27152 4380
rect 27152 4324 27156 4380
rect 27092 4320 27156 4324
rect 27172 4380 27236 4384
rect 27172 4324 27176 4380
rect 27176 4324 27232 4380
rect 27232 4324 27236 4380
rect 27172 4320 27236 4324
rect 27252 4380 27316 4384
rect 27252 4324 27256 4380
rect 27256 4324 27312 4380
rect 27312 4324 27316 4380
rect 27252 4320 27316 4324
rect 33012 4380 33076 4384
rect 33012 4324 33016 4380
rect 33016 4324 33072 4380
rect 33072 4324 33076 4380
rect 33012 4320 33076 4324
rect 33092 4380 33156 4384
rect 33092 4324 33096 4380
rect 33096 4324 33152 4380
rect 33152 4324 33156 4380
rect 33092 4320 33156 4324
rect 33172 4380 33236 4384
rect 33172 4324 33176 4380
rect 33176 4324 33232 4380
rect 33232 4324 33236 4380
rect 33172 4320 33236 4324
rect 33252 4380 33316 4384
rect 33252 4324 33256 4380
rect 33256 4324 33312 4380
rect 33312 4324 33316 4380
rect 33252 4320 33316 4324
rect 27660 4116 27724 4180
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 13952 3836 14016 3840
rect 13952 3780 13956 3836
rect 13956 3780 14012 3836
rect 14012 3780 14016 3836
rect 13952 3776 14016 3780
rect 14032 3836 14096 3840
rect 14032 3780 14036 3836
rect 14036 3780 14092 3836
rect 14092 3780 14096 3836
rect 14032 3776 14096 3780
rect 14112 3836 14176 3840
rect 14112 3780 14116 3836
rect 14116 3780 14172 3836
rect 14172 3780 14176 3836
rect 14112 3776 14176 3780
rect 14192 3836 14256 3840
rect 14192 3780 14196 3836
rect 14196 3780 14252 3836
rect 14252 3780 14256 3836
rect 14192 3776 14256 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 20192 3836 20256 3840
rect 20192 3780 20196 3836
rect 20196 3780 20252 3836
rect 20252 3780 20256 3836
rect 20192 3776 20256 3780
rect 25952 3836 26016 3840
rect 25952 3780 25956 3836
rect 25956 3780 26012 3836
rect 26012 3780 26016 3836
rect 25952 3776 26016 3780
rect 26032 3836 26096 3840
rect 26032 3780 26036 3836
rect 26036 3780 26092 3836
rect 26092 3780 26096 3836
rect 26032 3776 26096 3780
rect 26112 3836 26176 3840
rect 26112 3780 26116 3836
rect 26116 3780 26172 3836
rect 26172 3780 26176 3836
rect 26112 3776 26176 3780
rect 26192 3836 26256 3840
rect 26192 3780 26196 3836
rect 26196 3780 26252 3836
rect 26252 3780 26256 3836
rect 26192 3776 26256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 9172 3292 9236 3296
rect 9172 3236 9176 3292
rect 9176 3236 9232 3292
rect 9232 3236 9236 3292
rect 9172 3232 9236 3236
rect 9252 3292 9316 3296
rect 9252 3236 9256 3292
rect 9256 3236 9312 3292
rect 9312 3236 9316 3292
rect 9252 3232 9316 3236
rect 15012 3292 15076 3296
rect 15012 3236 15016 3292
rect 15016 3236 15072 3292
rect 15072 3236 15076 3292
rect 15012 3232 15076 3236
rect 15092 3292 15156 3296
rect 15092 3236 15096 3292
rect 15096 3236 15152 3292
rect 15152 3236 15156 3292
rect 15092 3232 15156 3236
rect 15172 3292 15236 3296
rect 15172 3236 15176 3292
rect 15176 3236 15232 3292
rect 15232 3236 15236 3292
rect 15172 3232 15236 3236
rect 15252 3292 15316 3296
rect 15252 3236 15256 3292
rect 15256 3236 15312 3292
rect 15312 3236 15316 3292
rect 15252 3232 15316 3236
rect 21012 3292 21076 3296
rect 21012 3236 21016 3292
rect 21016 3236 21072 3292
rect 21072 3236 21076 3292
rect 21012 3232 21076 3236
rect 21092 3292 21156 3296
rect 21092 3236 21096 3292
rect 21096 3236 21152 3292
rect 21152 3236 21156 3292
rect 21092 3232 21156 3236
rect 21172 3292 21236 3296
rect 21172 3236 21176 3292
rect 21176 3236 21232 3292
rect 21232 3236 21236 3292
rect 21172 3232 21236 3236
rect 21252 3292 21316 3296
rect 21252 3236 21256 3292
rect 21256 3236 21312 3292
rect 21312 3236 21316 3292
rect 21252 3232 21316 3236
rect 27012 3292 27076 3296
rect 27012 3236 27016 3292
rect 27016 3236 27072 3292
rect 27072 3236 27076 3292
rect 27012 3232 27076 3236
rect 27092 3292 27156 3296
rect 27092 3236 27096 3292
rect 27096 3236 27152 3292
rect 27152 3236 27156 3292
rect 27092 3232 27156 3236
rect 27172 3292 27236 3296
rect 27172 3236 27176 3292
rect 27176 3236 27232 3292
rect 27232 3236 27236 3292
rect 27172 3232 27236 3236
rect 27252 3292 27316 3296
rect 27252 3236 27256 3292
rect 27256 3236 27312 3292
rect 27312 3236 27316 3292
rect 27252 3232 27316 3236
rect 33012 3292 33076 3296
rect 33012 3236 33016 3292
rect 33016 3236 33072 3292
rect 33072 3236 33076 3292
rect 33012 3232 33076 3236
rect 33092 3292 33156 3296
rect 33092 3236 33096 3292
rect 33096 3236 33152 3292
rect 33152 3236 33156 3292
rect 33092 3232 33156 3236
rect 33172 3292 33236 3296
rect 33172 3236 33176 3292
rect 33176 3236 33232 3292
rect 33232 3236 33236 3292
rect 33172 3232 33236 3236
rect 33252 3292 33316 3296
rect 33252 3236 33256 3292
rect 33256 3236 33312 3292
rect 33312 3236 33316 3292
rect 33252 3232 33316 3236
rect 25636 2892 25700 2956
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 13952 2748 14016 2752
rect 13952 2692 13956 2748
rect 13956 2692 14012 2748
rect 14012 2692 14016 2748
rect 13952 2688 14016 2692
rect 14032 2748 14096 2752
rect 14032 2692 14036 2748
rect 14036 2692 14092 2748
rect 14092 2692 14096 2748
rect 14032 2688 14096 2692
rect 14112 2748 14176 2752
rect 14112 2692 14116 2748
rect 14116 2692 14172 2748
rect 14172 2692 14176 2748
rect 14112 2688 14176 2692
rect 14192 2748 14256 2752
rect 14192 2692 14196 2748
rect 14196 2692 14252 2748
rect 14252 2692 14256 2748
rect 14192 2688 14256 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 20192 2748 20256 2752
rect 20192 2692 20196 2748
rect 20196 2692 20252 2748
rect 20252 2692 20256 2748
rect 20192 2688 20256 2692
rect 25952 2748 26016 2752
rect 25952 2692 25956 2748
rect 25956 2692 26012 2748
rect 26012 2692 26016 2748
rect 25952 2688 26016 2692
rect 26032 2748 26096 2752
rect 26032 2692 26036 2748
rect 26036 2692 26092 2748
rect 26092 2692 26096 2748
rect 26032 2688 26096 2692
rect 26112 2748 26176 2752
rect 26112 2692 26116 2748
rect 26116 2692 26172 2748
rect 26172 2692 26176 2748
rect 26112 2688 26176 2692
rect 26192 2748 26256 2752
rect 26192 2692 26196 2748
rect 26196 2692 26252 2748
rect 26252 2692 26256 2748
rect 26192 2688 26256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 26740 2484 26804 2548
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 9172 2204 9236 2208
rect 9172 2148 9176 2204
rect 9176 2148 9232 2204
rect 9232 2148 9236 2204
rect 9172 2144 9236 2148
rect 9252 2204 9316 2208
rect 9252 2148 9256 2204
rect 9256 2148 9312 2204
rect 9312 2148 9316 2204
rect 9252 2144 9316 2148
rect 15012 2204 15076 2208
rect 15012 2148 15016 2204
rect 15016 2148 15072 2204
rect 15072 2148 15076 2204
rect 15012 2144 15076 2148
rect 15092 2204 15156 2208
rect 15092 2148 15096 2204
rect 15096 2148 15152 2204
rect 15152 2148 15156 2204
rect 15092 2144 15156 2148
rect 15172 2204 15236 2208
rect 15172 2148 15176 2204
rect 15176 2148 15232 2204
rect 15232 2148 15236 2204
rect 15172 2144 15236 2148
rect 15252 2204 15316 2208
rect 15252 2148 15256 2204
rect 15256 2148 15312 2204
rect 15312 2148 15316 2204
rect 15252 2144 15316 2148
rect 21012 2204 21076 2208
rect 21012 2148 21016 2204
rect 21016 2148 21072 2204
rect 21072 2148 21076 2204
rect 21012 2144 21076 2148
rect 21092 2204 21156 2208
rect 21092 2148 21096 2204
rect 21096 2148 21152 2204
rect 21152 2148 21156 2204
rect 21092 2144 21156 2148
rect 21172 2204 21236 2208
rect 21172 2148 21176 2204
rect 21176 2148 21232 2204
rect 21232 2148 21236 2204
rect 21172 2144 21236 2148
rect 21252 2204 21316 2208
rect 21252 2148 21256 2204
rect 21256 2148 21312 2204
rect 21312 2148 21316 2204
rect 21252 2144 21316 2148
rect 27012 2204 27076 2208
rect 27012 2148 27016 2204
rect 27016 2148 27072 2204
rect 27072 2148 27076 2204
rect 27012 2144 27076 2148
rect 27092 2204 27156 2208
rect 27092 2148 27096 2204
rect 27096 2148 27152 2204
rect 27152 2148 27156 2204
rect 27092 2144 27156 2148
rect 27172 2204 27236 2208
rect 27172 2148 27176 2204
rect 27176 2148 27232 2204
rect 27232 2148 27236 2204
rect 27172 2144 27236 2148
rect 27252 2204 27316 2208
rect 27252 2148 27256 2204
rect 27256 2148 27312 2204
rect 27312 2148 27316 2204
rect 27252 2144 27316 2148
rect 33012 2204 33076 2208
rect 33012 2148 33016 2204
rect 33016 2148 33072 2204
rect 33072 2148 33076 2204
rect 33012 2144 33076 2148
rect 33092 2204 33156 2208
rect 33092 2148 33096 2204
rect 33096 2148 33152 2204
rect 33152 2148 33156 2204
rect 33092 2144 33156 2148
rect 33172 2204 33236 2208
rect 33172 2148 33176 2204
rect 33176 2148 33232 2204
rect 33232 2148 33236 2204
rect 33172 2144 33236 2148
rect 33252 2204 33316 2208
rect 33252 2148 33256 2204
rect 33256 2148 33312 2204
rect 33312 2148 33316 2204
rect 33252 2144 33316 2148
rect 25636 580 25700 644
rect 28212 444 28276 508
rect 27660 172 27724 236
rect 25084 96 25148 100
rect 25084 40 25134 96
rect 25134 40 25148 96
rect 25084 36 25148 40
<< metal4 >>
rect 1944 8192 2264 11152
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 0 2264 2688
rect 3004 8736 3324 11152
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 0 3324 2144
rect 7944 8192 8264 11152
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 7944 6016 8264 7040
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 4928 8264 5952
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 2752 8264 3776
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 7944 0 8264 2688
rect 9004 8736 9324 11152
rect 9004 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9324 8736
rect 9004 7648 9324 8672
rect 9004 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9324 7648
rect 9004 6560 9324 7584
rect 9004 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9324 6560
rect 9004 5472 9324 6496
rect 9004 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9324 5472
rect 9004 4384 9324 5408
rect 9004 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9324 4384
rect 9004 3296 9324 4320
rect 9004 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9324 3296
rect 9004 2208 9324 3232
rect 9004 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9324 2208
rect 9004 0 9324 2144
rect 13944 8192 14264 11152
rect 13944 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14264 8192
rect 13944 7104 14264 8128
rect 13944 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14264 7104
rect 13944 6016 14264 7040
rect 13944 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14264 6016
rect 13944 4928 14264 5952
rect 13944 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14264 4928
rect 13944 3840 14264 4864
rect 13944 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14264 3840
rect 13944 2752 14264 3776
rect 13944 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14264 2752
rect 13944 0 14264 2688
rect 15004 8736 15324 11152
rect 15004 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15324 8736
rect 15004 7648 15324 8672
rect 15004 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15324 7648
rect 15004 6560 15324 7584
rect 15004 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15324 6560
rect 15004 5472 15324 6496
rect 15004 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15324 5472
rect 15004 4384 15324 5408
rect 15004 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15324 4384
rect 15004 3296 15324 4320
rect 15004 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15324 3296
rect 15004 2208 15324 3232
rect 15004 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15324 2208
rect 15004 0 15324 2144
rect 19944 8192 20264 11152
rect 19944 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20264 8192
rect 19944 7104 20264 8128
rect 19944 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20264 7104
rect 19944 6016 20264 7040
rect 19944 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20264 6016
rect 19944 4928 20264 5952
rect 19944 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20264 4928
rect 19944 3840 20264 4864
rect 19944 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20264 3840
rect 19944 2752 20264 3776
rect 19944 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20264 2752
rect 19944 0 20264 2688
rect 21004 8736 21324 11152
rect 21004 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21324 8736
rect 21004 7648 21324 8672
rect 21004 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21324 7648
rect 21004 6560 21324 7584
rect 21004 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21324 6560
rect 21004 5472 21324 6496
rect 25944 8192 26264 11152
rect 25944 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26264 8192
rect 25944 7104 26264 8128
rect 25944 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26264 7104
rect 25944 6016 26264 7040
rect 25944 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26264 6016
rect 25083 5812 25149 5813
rect 25083 5748 25084 5812
rect 25148 5748 25149 5812
rect 25083 5747 25149 5748
rect 21004 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21324 5472
rect 21004 4384 21324 5408
rect 21004 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21324 4384
rect 21004 3296 21324 4320
rect 21004 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21324 3296
rect 21004 2208 21324 3232
rect 21004 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21324 2208
rect 21004 0 21324 2144
rect 25086 101 25146 5747
rect 25944 4928 26264 5952
rect 25944 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26264 4928
rect 25944 3840 26264 4864
rect 27004 8736 27324 11152
rect 27004 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27324 8736
rect 27004 7648 27324 8672
rect 27004 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27324 7648
rect 27004 6560 27324 7584
rect 27004 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27324 6560
rect 27004 5472 27324 6496
rect 27004 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27324 5472
rect 26739 4724 26805 4725
rect 26739 4660 26740 4724
rect 26804 4660 26805 4724
rect 26739 4659 26805 4660
rect 25944 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26264 3840
rect 25635 2956 25701 2957
rect 25635 2892 25636 2956
rect 25700 2892 25701 2956
rect 25635 2891 25701 2892
rect 25638 645 25698 2891
rect 25944 2752 26264 3776
rect 25944 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26264 2752
rect 25635 644 25701 645
rect 25635 580 25636 644
rect 25700 580 25701 644
rect 25635 579 25701 580
rect 25083 100 25149 101
rect 25083 36 25084 100
rect 25148 36 25149 100
rect 25083 35 25149 36
rect 25944 0 26264 2688
rect 26742 2549 26802 4659
rect 27004 4384 27324 5408
rect 31944 8192 32264 11152
rect 31944 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32264 8192
rect 31944 7104 32264 8128
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 28211 4588 28277 4589
rect 28211 4524 28212 4588
rect 28276 4524 28277 4588
rect 28211 4523 28277 4524
rect 27004 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27324 4384
rect 27004 3296 27324 4320
rect 27659 4180 27725 4181
rect 27659 4116 27660 4180
rect 27724 4116 27725 4180
rect 27659 4115 27725 4116
rect 27004 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27324 3296
rect 26739 2548 26805 2549
rect 26739 2484 26740 2548
rect 26804 2484 26805 2548
rect 26739 2483 26805 2484
rect 27004 2208 27324 3232
rect 27004 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27324 2208
rect 27004 0 27324 2144
rect 27662 237 27722 4115
rect 28214 509 28274 4523
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 2752 32264 3776
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 28211 508 28277 509
rect 28211 444 28212 508
rect 28276 444 28277 508
rect 28211 443 28277 444
rect 27659 236 27725 237
rect 27659 172 27660 236
rect 27724 172 27725 236
rect 27659 171 27725 172
rect 31944 0 32264 2688
rect 33004 8736 33324 11152
rect 33004 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33324 8736
rect 33004 7648 33324 8672
rect 33004 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33324 7648
rect 33004 6560 33324 7584
rect 33004 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33324 6560
rect 33004 5472 33324 6496
rect 33004 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33324 5472
rect 33004 4384 33324 5408
rect 33004 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33324 4384
rect 33004 3296 33324 4320
rect 33004 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33324 3296
rect 33004 2208 33324 3232
rect 33004 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33324 2208
rect 33004 0 33324 2144
use sky130_fd_sc_hd__buf_1  _000_
timestamp -3599
transform 1 0 17940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _001_
timestamp -3599
transform 1 0 20976 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _002_
timestamp -3599
transform 1 0 21528 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _003_
timestamp -3599
transform 1 0 21804 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _004_
timestamp -3599
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _005_
timestamp -3599
transform -1 0 24932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _006_
timestamp -3599
transform -1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _007_
timestamp -3599
transform -1 0 24196 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _008_
timestamp -3599
transform -1 0 25208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _009_
timestamp -3599
transform 1 0 21252 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _010_
timestamp -3599
transform 1 0 23920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _011_
timestamp -3599
transform 1 0 24196 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _012_
timestamp -3599
transform -1 0 24748 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _013_
timestamp -3599
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _014_
timestamp -3599
transform 1 0 17756 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _015_
timestamp -3599
transform 1 0 18032 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _016_
timestamp -3599
transform 1 0 19780 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _017_
timestamp -3599
transform 1 0 22448 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _018_
timestamp -3599
transform 1 0 16744 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _019_
timestamp -3599
transform 1 0 18676 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _020_
timestamp -3599
transform 1 0 16376 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _021_
timestamp -3599
transform 1 0 15732 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _022_
timestamp -3599
transform 1 0 21436 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _023_
timestamp -3599
transform 1 0 15456 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _024_
timestamp -3599
transform 1 0 18952 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _025_
timestamp -3599
transform 1 0 18124 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _026_
timestamp -3599
transform 1 0 20240 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _027_
timestamp -3599
transform 1 0 17204 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _028_
timestamp -3599
transform 1 0 17480 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _029_
timestamp -3599
transform 1 0 15364 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _030_
timestamp -3599
transform 1 0 17020 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _031_
timestamp -3599
transform 1 0 21160 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _032_
timestamp -3599
transform 1 0 9292 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _033_
timestamp -3599
transform 1 0 12144 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _034_
timestamp -3599
transform 1 0 14812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _035_
timestamp -3599
transform 1 0 14168 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _036_
timestamp -3599
transform -1 0 25024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _037_
timestamp -3599
transform -1 0 28520 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _038_
timestamp -3599
transform -1 0 28796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _039_
timestamp -3599
transform -1 0 26312 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _040_
timestamp -3599
transform 1 0 25116 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _041_
timestamp -3599
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _042_
timestamp -3599
transform 1 0 25300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _043_
timestamp -3599
transform 1 0 27692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _044_
timestamp -3599
transform 1 0 29440 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp -3599
transform 1 0 30912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp -3599
transform -1 0 24932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _047_
timestamp -3599
transform 1 0 27968 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp -3599
transform 1 0 28704 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp -3599
transform 1 0 29716 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _050_
timestamp -3599
transform -1 0 31096 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _051_
timestamp -3599
transform -1 0 28980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _052_
timestamp -3599
transform 1 0 2944 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _053_
timestamp -3599
transform 1 0 3220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _054_
timestamp -3599
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _055_
timestamp -3599
transform 1 0 2944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _056_
timestamp -3599
transform 1 0 2484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _057_
timestamp -3599
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _058_
timestamp -3599
transform 1 0 1932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _059_
timestamp -3599
transform 1 0 2300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _060_
timestamp -3599
transform 1 0 3404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _061_
timestamp -3599
transform 1 0 3680 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _062_
timestamp -3599
transform 1 0 4232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _063_
timestamp -3599
transform 1 0 4600 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _064_
timestamp -3599
transform 1 0 6532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _065_
timestamp -3599
transform 1 0 7176 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _066_
timestamp -3599
transform 1 0 7176 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _067_
timestamp -3599
transform 1 0 6808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _068_
timestamp -3599
transform 1 0 7084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _069_
timestamp -3599
transform 1 0 7912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _070_
timestamp -3599
transform 1 0 7636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _071_
timestamp -3599
transform 1 0 7360 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp -3599
transform -1 0 15272 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp -3599
transform -1 0 14996 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp -3599
transform -1 0 11040 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp -3599
transform -1 0 11316 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp -3599
transform -1 0 11592 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp -3599
transform -1 0 11868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp -3599
transform -1 0 12144 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp -3599
transform -1 0 12512 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp -3599
transform -1 0 12788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp -3599
transform -1 0 13616 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp -3599
transform -1 0 13340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp -3599
transform -1 0 13892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp -3599
transform -1 0 14260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp -3599
transform -1 0 14720 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp -3599
transform -1 0 15640 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp -3599
transform -1 0 15364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp -3599
transform 1 0 29348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp -3599
transform 1 0 28244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp -3599
transform 1 0 28704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp -3599
transform 1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp -3599
transform 1 0 27968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp -3599
transform 1 0 28612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp -3599
transform 1 0 27692 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp -3599
transform 1 0 27600 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp -3599
transform 1 0 28428 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp -3599
transform 1 0 28060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp -3599
transform 1 0 27784 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp -3599
transform 1 0 27508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp -3599
transform 1 0 27232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp -3599
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp -3599
transform 1 0 26680 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp -3599
transform 1 0 26404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp -3599
transform -1 0 11316 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform -1 0 17940 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform 1 0 17572 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform 1 0 22264 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform -1 0 16560 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform -1 0 18676 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform -1 0 20976 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform 1 0 16192 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform -1 0 16192 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp -3599
transform 1 0 20700 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp -3599
transform 1 0 15272 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp -3599
transform -1 0 19412 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp -3599
transform 1 0 17020 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp -3599
transform -1 0 17940 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp -3599
transform -1 0 15364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp -3599
transform -1 0 22264 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp -3599
transform -1 0 17480 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp -3599
transform -1 0 22448 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp -3599
transform -1 0 19688 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp -3599
transform -1 0 25392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp -3599
transform -1 0 23920 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp -3599
transform -1 0 23736 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp -3599
transform -1 0 25576 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp -3599
transform 1 0 20608 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp -3599
transform -1 0 9292 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp -3599
transform -1 0 14812 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp -3599
transform 1 0 28428 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp -3599
transform -1 0 27968 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp -3599
transform -1 0 29348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp -3599
transform -1 0 28152 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp -3599
transform -1 0 28704 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp -3599
transform 1 0 27600 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp -3599
transform 1 0 27416 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp -3599
transform 1 0 20976 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp -3599
transform -1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp -3599
transform -1 0 10948 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3
timestamp -3599
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6
timestamp -3599
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9
timestamp -3599
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12
timestamp -3599
transform 1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15
timestamp -3599
transform 1 0 2484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18
timestamp -3599
transform 1 0 2760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21
timestamp -3599
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24
timestamp -3599
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29
timestamp -3599
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp -3599
transform 1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35
timestamp -3599
transform 1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38
timestamp -3599
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41
timestamp -3599
transform 1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44
timestamp -3599
transform 1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47
timestamp -3599
transform 1 0 5428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50
timestamp -3599
transform 1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -3599
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp -3599
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60
timestamp -3599
transform 1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63
timestamp -3599
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66
timestamp -3599
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69
timestamp -3599
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72
timestamp -3599
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75
timestamp -3599
transform 1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_78
timestamp -3599
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -3599
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85
timestamp -3599
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_88
timestamp -3599
transform 1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_91
timestamp -3599
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_94
timestamp -3599
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_97
timestamp -3599
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100
timestamp -3599
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_103
timestamp -3599
transform 1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_106
timestamp -3599
transform 1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -3599
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp -3599
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_116
timestamp -3599
transform 1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119
timestamp -3599
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_122
timestamp -3599
transform 1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_125
timestamp -3599
transform 1 0 12604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_128
timestamp -3599
transform 1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_131
timestamp -3599
transform 1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_134
timestamp -3599
transform 1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp -3599
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141
timestamp -3599
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_144
timestamp -3599
transform 1 0 14352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_147
timestamp -3599
transform 1 0 14628 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp -3599
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp -3599
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp -3599
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_273
timestamp -3599
transform 1 0 26220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_276
timestamp -3599
transform 1 0 26496 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp -3599
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_281
timestamp -3599
transform 1 0 26956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_284
timestamp -3599
transform 1 0 27232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_287
timestamp -3599
transform 1 0 27508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_290
timestamp -3599
transform 1 0 27784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_293
timestamp -3599
transform 1 0 28060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_296
timestamp -3599
transform 1 0 28336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_299
timestamp -3599
transform 1 0 28612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_302
timestamp -3599
transform 1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp -3599
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_309
timestamp -3599
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_312
timestamp -3599
transform 1 0 29808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_315
timestamp -3599
transform 1 0 30084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_318
timestamp -3599
transform 1 0 30360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_321
timestamp -3599
transform 1 0 30636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp -3599
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp -3599
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_6
timestamp -3599
transform 1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_9
timestamp -3599
transform 1 0 1932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_12
timestamp -3599
transform 1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_15
timestamp -3599
transform 1 0 2484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_18
timestamp -3599
transform 1 0 2760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_21
timestamp -3599
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_24
timestamp -3599
transform 1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_27
timestamp -3599
transform 1 0 3588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_30
timestamp -3599
transform 1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_33
timestamp -3599
transform 1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_36
timestamp -3599
transform 1 0 4416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_39
timestamp -3599
transform 1 0 4692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_42
timestamp -3599
transform 1 0 4968 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_45
timestamp -3599
transform 1 0 5244 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_48
timestamp -3599
transform 1 0 5520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_51
timestamp -3599
transform 1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp -3599
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp -3599
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_60
timestamp -3599
transform 1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_63
timestamp -3599
transform 1 0 6900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_66
timestamp -3599
transform 1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_69
timestamp -3599
transform 1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_72
timestamp -3599
transform 1 0 7728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_75
timestamp -3599
transform 1 0 8004 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_78
timestamp -3599
transform 1 0 8280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_81
timestamp -3599
transform 1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_84
timestamp -3599
transform 1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_87
timestamp -3599
transform 1 0 9108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_90
timestamp -3599
transform 1 0 9384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_93
timestamp -3599
transform 1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_96
timestamp -3599
transform 1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_99
timestamp -3599
transform 1 0 10212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_102
timestamp -3599
transform 1 0 10488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_105
timestamp -3599
transform 1 0 10764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_108
timestamp -3599
transform 1 0 11040 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp -3599
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp -3599
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_116
timestamp -3599
transform 1 0 11776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_119
timestamp -3599
transform 1 0 12052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_122
timestamp -3599
transform 1 0 12328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_125
timestamp -3599
transform 1 0 12604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_128
timestamp -3599
transform 1 0 12880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_131
timestamp -3599
transform 1 0 13156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_134
timestamp -3599
transform 1 0 13432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_137
timestamp -3599
transform 1 0 13708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_140
timestamp -3599
transform 1 0 13984 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_143
timestamp -3599
transform 1 0 14260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_146
timestamp -3599
transform 1 0 14536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_149
timestamp -3599
transform 1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_152
timestamp -3599
transform 1 0 15088 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_155
timestamp -3599
transform 1 0 15364 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_169
timestamp -3599
transform 1 0 16652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_182
timestamp -3599
transform 1 0 17848 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_185
timestamp -3599
transform 1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_188
timestamp -3599
transform 1 0 18400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_191
timestamp -3599
transform 1 0 18676 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp -3599
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_269
timestamp -3599
transform 1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_272
timestamp -3599
transform 1 0 26128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_275
timestamp -3599
transform 1 0 26404 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp -3599
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_281
timestamp -3599
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_284
timestamp -3599
transform 1 0 27232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_287
timestamp -3599
transform 1 0 27508 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_291
timestamp -3599
transform 1 0 27876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_294
timestamp -3599
transform 1 0 28152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_297
timestamp -3599
transform 1 0 28428 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_300
timestamp -3599
transform 1 0 28704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_303
timestamp -3599
transform 1 0 28980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_306
timestamp -3599
transform 1 0 29256 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_309
timestamp -3599
transform 1 0 29532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_312
timestamp -3599
transform 1 0 29808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_315
timestamp -3599
transform 1 0 30084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_318
timestamp -3599
transform 1 0 30360 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_321
timestamp -3599
transform 1 0 30636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_324
timestamp -3599
transform 1 0 30912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_327
timestamp -3599
transform 1 0 31188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_330
timestamp -3599
transform 1 0 31464 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp -3599
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp -3599
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_6
timestamp -3599
transform 1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_9
timestamp -3599
transform 1 0 1932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_12
timestamp -3599
transform 1 0 2208 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_16
timestamp -3599
transform 1 0 2576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_19
timestamp -3599
transform 1 0 2852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_22
timestamp -3599
transform 1 0 3128 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_25
timestamp -3599
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_29
timestamp -3599
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_32
timestamp -3599
transform 1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_35
timestamp -3599
transform 1 0 4324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_38
timestamp -3599
transform 1 0 4600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_41
timestamp -3599
transform 1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_44
timestamp -3599
transform 1 0 5152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_47
timestamp -3599
transform 1 0 5428 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_50
timestamp -3599
transform 1 0 5704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_53
timestamp -3599
transform 1 0 5980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_56
timestamp -3599
transform 1 0 6256 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_59
timestamp -3599
transform 1 0 6532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_62
timestamp -3599
transform 1 0 6808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_65
timestamp -3599
transform 1 0 7084 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_69
timestamp -3599
transform 1 0 7452 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_72
timestamp -3599
transform 1 0 7728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_75
timestamp -3599
transform 1 0 8004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_78
timestamp -3599
transform 1 0 8280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp -3599
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_85
timestamp -3599
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_88
timestamp -3599
transform 1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_91
timestamp -3599
transform 1 0 9476 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_94
timestamp -3599
transform 1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_97
timestamp -3599
transform 1 0 10028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_100
timestamp -3599
transform 1 0 10304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_103
timestamp -3599
transform 1 0 10580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_106
timestamp -3599
transform 1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_109
timestamp -3599
transform 1 0 11132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_112
timestamp -3599
transform 1 0 11408 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_115
timestamp -3599
transform 1 0 11684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_118
timestamp -3599
transform 1 0 11960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_121
timestamp -3599
transform 1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_124
timestamp -3599
transform 1 0 12512 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_127
timestamp -3599
transform 1 0 12788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_130
timestamp -3599
transform 1 0 13064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_133
timestamp -3599
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_136
timestamp -3599
transform 1 0 13616 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp -3599
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_141
timestamp -3599
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_144
timestamp -3599
transform 1 0 14352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_147
timestamp -3599
transform 1 0 14628 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_150
timestamp -3599
transform 1 0 14904 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_153
timestamp -3599
transform 1 0 15180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_156
timestamp -3599
transform 1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_159
timestamp -3599
transform 1 0 15732 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_162
timestamp -3599
transform 1 0 16008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_165
timestamp -3599
transform 1 0 16284 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_168
timestamp -3599
transform 1 0 16560 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_171
timestamp -3599
transform 1 0 16836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_174
timestamp -3599
transform 1 0 17112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_177
timestamp -3599
transform 1 0 17388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_180
timestamp -3599
transform 1 0 17664 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_186
timestamp -3599
transform 1 0 18216 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_189
timestamp -3599
transform 1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_192
timestamp -3599
transform 1 0 18768 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp -3599
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_202
timestamp -3599
transform 1 0 19688 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_205
timestamp -3599
transform 1 0 19964 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_208
timestamp -3599
transform 1 0 20240 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_211
timestamp -3599
transform 1 0 20516 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_232
timestamp -3599
transform 1 0 22448 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_235
timestamp -3599
transform 1 0 22724 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_238
timestamp -3599
transform 1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_241
timestamp -3599
transform 1 0 23276 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp -3599
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_266
timestamp -3599
transform 1 0 25576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_269
timestamp -3599
transform 1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_272
timestamp -3599
transform 1 0 26128 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_281
timestamp -3599
transform 1 0 26956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_300
timestamp -3599
transform 1 0 28704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_303
timestamp -3599
transform 1 0 28980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp -3599
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_309
timestamp -3599
transform 1 0 29532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_312
timestamp -3599
transform 1 0 29808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_315
timestamp -3599
transform 1 0 30084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_318
timestamp -3599
transform 1 0 30360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_321
timestamp -3599
transform 1 0 30636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_324
timestamp -3599
transform 1 0 30912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_327
timestamp -3599
transform 1 0 31188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_330
timestamp -3599
transform 1 0 31464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_333
timestamp -3599
transform 1 0 31740 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_336
timestamp -3599
transform 1 0 32016 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp -3599
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_6
timestamp -3599
transform 1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_18
timestamp -3599
transform 1 0 2760 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_23
timestamp -3599
transform 1 0 3220 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_31
timestamp -3599
transform 1 0 3956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_37
timestamp -3599
transform 1 0 4508 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_41
timestamp -3599
transform 1 0 4876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_44
timestamp -3599
transform 1 0 5152 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_47
timestamp -3599
transform 1 0 5428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_50
timestamp -3599
transform 1 0 5704 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp -3599
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp -3599
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_77
timestamp -3599
transform 1 0 8188 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_80
timestamp -3599
transform 1 0 8464 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_83
timestamp -3599
transform 1 0 8740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_86
timestamp -3599
transform 1 0 9016 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_89
timestamp -3599
transform 1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_92
timestamp -3599
transform 1 0 9568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_95
timestamp -3599
transform 1 0 9844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_98
timestamp -3599
transform 1 0 10120 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_101
timestamp -3599
transform 1 0 10396 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_104
timestamp -3599
transform 1 0 10672 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_107
timestamp -3599
transform 1 0 10948 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp -3599
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_113
timestamp -3599
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_116
timestamp -3599
transform 1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp -3599
transform 1 0 12052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_122
timestamp -3599
transform 1 0 12328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_125
timestamp -3599
transform 1 0 12604 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_128
timestamp -3599
transform 1 0 12880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_131
timestamp -3599
transform 1 0 13156 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_134
timestamp -3599
transform 1 0 13432 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_137
timestamp -3599
transform 1 0 13708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_143
timestamp -3599
transform 1 0 14260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_148
timestamp -3599
transform 1 0 14720 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_151
timestamp -3599
transform 1 0 14996 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_158
timestamp -3599
transform 1 0 15640 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_161
timestamp -3599
transform 1 0 15916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_164
timestamp -3599
transform 1 0 16192 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp -3599
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_169
timestamp -3599
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_172
timestamp -3599
transform 1 0 16928 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_175
timestamp -3599
transform 1 0 17204 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_178
timestamp -3599
transform 1 0 17480 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_181
timestamp -3599
transform 1 0 17756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_184
timestamp -3599
transform 1 0 18032 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_187
timestamp -3599
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_190
timestamp -3599
transform 1 0 18584 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_193
timestamp -3599
transform 1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_196
timestamp -3599
transform 1 0 19136 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_199
timestamp -3599
transform 1 0 19412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_202
timestamp -3599
transform 1 0 19688 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_205
timestamp -3599
transform 1 0 19964 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_208
timestamp -3599
transform 1 0 20240 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_211
timestamp -3599
transform 1 0 20516 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_214
timestamp -3599
transform 1 0 20792 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_217
timestamp -3599
transform 1 0 21068 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_220
timestamp -3599
transform 1 0 21344 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp -3599
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp -3599
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_228
timestamp -3599
transform 1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_231
timestamp -3599
transform 1 0 22356 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_234
timestamp -3599
transform 1 0 22632 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_237
timestamp -3599
transform 1 0 22908 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_240
timestamp -3599
transform 1 0 23184 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_243
timestamp -3599
transform 1 0 23460 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_246
timestamp -3599
transform 1 0 23736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_249
timestamp -3599
transform 1 0 24012 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_252
timestamp -3599
transform 1 0 24288 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_255
timestamp -3599
transform 1 0 24564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_258
timestamp -3599
transform 1 0 24840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_261
timestamp -3599
transform 1 0 25116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_264
timestamp -3599
transform 1 0 25392 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_267
timestamp -3599
transform 1 0 25668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_270
timestamp -3599
transform 1 0 25944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_273
timestamp -3599
transform 1 0 26220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_276
timestamp -3599
transform 1 0 26496 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp -3599
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_284
timestamp -3599
transform 1 0 27232 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_296
timestamp -3599
transform 1 0 28336 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_310
timestamp -3599
transform 1 0 29624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_313
timestamp -3599
transform 1 0 29900 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_316
timestamp -3599
transform 1 0 30176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_319
timestamp -3599
transform 1 0 30452 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_322
timestamp -3599
transform 1 0 30728 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_325
timestamp -3599
transform 1 0 31004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_328
timestamp -3599
transform 1 0 31280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_331
timestamp -3599
transform 1 0 31556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp -3599
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp -3599
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp -3599
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_6
timestamp -3599
transform 1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_9
timestamp -3599
transform 1 0 1932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_12
timestamp -3599
transform 1 0 2208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_15
timestamp -3599
transform 1 0 2484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_18
timestamp -3599
transform 1 0 2760 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp -3599
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_32
timestamp -3599
transform 1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_35
timestamp -3599
transform 1 0 4324 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_38
timestamp -3599
transform 1 0 4600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_41
timestamp -3599
transform 1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_44
timestamp -3599
transform 1 0 5152 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_47
timestamp -3599
transform 1 0 5428 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_50
timestamp -3599
transform 1 0 5704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_53
timestamp -3599
transform 1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_56
timestamp -3599
transform 1 0 6256 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_59
timestamp -3599
transform 1 0 6532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_62
timestamp -3599
transform 1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_65
timestamp -3599
transform 1 0 7084 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_69
timestamp -3599
transform 1 0 7452 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_72
timestamp -3599
transform 1 0 7728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_75
timestamp -3599
transform 1 0 8004 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_78
timestamp -3599
transform 1 0 8280 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp -3599
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_85
timestamp -3599
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_88
timestamp -3599
transform 1 0 9200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_91
timestamp -3599
transform 1 0 9476 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_94
timestamp -3599
transform 1 0 9752 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_97
timestamp -3599
transform 1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_100
timestamp -3599
transform 1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_103
timestamp -3599
transform 1 0 10580 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_120
timestamp -3599
transform 1 0 12144 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_127
timestamp -3599
transform 1 0 12788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp -3599
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_141
timestamp -3599
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_144
timestamp -3599
transform 1 0 14352 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_147
timestamp -3599
transform 1 0 14628 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_169
timestamp -3599
transform 1 0 16652 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_172
timestamp -3599
transform 1 0 16928 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_175
timestamp -3599
transform 1 0 17204 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_178
timestamp -3599
transform 1 0 17480 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_181
timestamp -3599
transform 1 0 17756 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_184
timestamp -3599
transform 1 0 18032 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_187
timestamp -3599
transform 1 0 18308 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_190
timestamp -3599
transform 1 0 18584 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp -3599
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp -3599
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_200
timestamp -3599
transform 1 0 19504 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_203
timestamp -3599
transform 1 0 19780 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_206
timestamp -3599
transform 1 0 20056 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_209
timestamp -3599
transform 1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_212
timestamp -3599
transform 1 0 20608 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_215
timestamp -3599
transform 1 0 20884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_218
timestamp -3599
transform 1 0 21160 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_221
timestamp -3599
transform 1 0 21436 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_224
timestamp -3599
transform 1 0 21712 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_227
timestamp -3599
transform 1 0 21988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_230
timestamp -3599
transform 1 0 22264 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_233
timestamp -3599
transform 1 0 22540 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_236
timestamp -3599
transform 1 0 22816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_239
timestamp -3599
transform 1 0 23092 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_242
timestamp -3599
transform 1 0 23368 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_245
timestamp -3599
transform 1 0 23644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_248
timestamp -3599
transform 1 0 23920 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp -3599
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_253
timestamp -3599
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_256
timestamp -3599
transform 1 0 24656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_259
timestamp -3599
transform 1 0 24932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_262
timestamp -3599
transform 1 0 25208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_265
timestamp -3599
transform 1 0 25484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_268
timestamp -3599
transform 1 0 25760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_271
timestamp -3599
transform 1 0 26036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_274
timestamp -3599
transform 1 0 26312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_277
timestamp -3599
transform 1 0 26588 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_280
timestamp -3599
transform 1 0 26864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_283
timestamp -3599
transform 1 0 27140 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_286
timestamp -3599
transform 1 0 27416 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_294
timestamp -3599
transform 1 0 28152 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_303
timestamp -3599
transform 1 0 28980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp -3599
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_309
timestamp -3599
transform 1 0 29532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_312
timestamp -3599
transform 1 0 29808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_315
timestamp -3599
transform 1 0 30084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_318
timestamp -3599
transform 1 0 30360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_321
timestamp -3599
transform 1 0 30636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_324
timestamp -3599
transform 1 0 30912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_327
timestamp -3599
transform 1 0 31188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_330
timestamp -3599
transform 1 0 31464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_333
timestamp -3599
transform 1 0 31740 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_336
timestamp -3599
transform 1 0 32016 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp -3599
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_6
timestamp -3599
transform 1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_9
timestamp -3599
transform 1 0 1932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_12
timestamp -3599
transform 1 0 2208 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_15
timestamp -3599
transform 1 0 2484 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_18
timestamp -3599
transform 1 0 2760 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_21
timestamp -3599
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_24
timestamp -3599
transform 1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_27
timestamp -3599
transform 1 0 3588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_30
timestamp -3599
transform 1 0 3864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_33
timestamp -3599
transform 1 0 4140 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_36
timestamp -3599
transform 1 0 4416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_39
timestamp -3599
transform 1 0 4692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_42
timestamp -3599
transform 1 0 4968 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_45
timestamp -3599
transform 1 0 5244 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_48
timestamp -3599
transform 1 0 5520 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_51
timestamp -3599
transform 1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp -3599
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_57
timestamp -3599
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_60
timestamp -3599
transform 1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_63
timestamp -3599
transform 1 0 6900 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_66
timestamp -3599
transform 1 0 7176 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_69
timestamp -3599
transform 1 0 7452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_72
timestamp -3599
transform 1 0 7728 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_75
timestamp -3599
transform 1 0 8004 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_78
timestamp -3599
transform 1 0 8280 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_81
timestamp -3599
transform 1 0 8556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_84
timestamp -3599
transform 1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_87
timestamp -3599
transform 1 0 9108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_90
timestamp -3599
transform 1 0 9384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_93
timestamp -3599
transform 1 0 9660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_96
timestamp -3599
transform 1 0 9936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_99
timestamp -3599
transform 1 0 10212 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_102
timestamp -3599
transform 1 0 10488 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_105
timestamp -3599
transform 1 0 10764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_108
timestamp -3599
transform 1 0 11040 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp -3599
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_113
timestamp -3599
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_116
timestamp -3599
transform 1 0 11776 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_119
timestamp -3599
transform 1 0 12052 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_122
timestamp -3599
transform 1 0 12328 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_125
timestamp -3599
transform 1 0 12604 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_128
timestamp -3599
transform 1 0 12880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_131
timestamp -3599
transform 1 0 13156 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_134
timestamp -3599
transform 1 0 13432 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_137
timestamp -3599
transform 1 0 13708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_140
timestamp -3599
transform 1 0 13984 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_143
timestamp -3599
transform 1 0 14260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_146
timestamp -3599
transform 1 0 14536 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_149
timestamp -3599
transform 1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_152
timestamp -3599
transform 1 0 15088 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_158
timestamp -3599
transform 1 0 15640 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_161
timestamp -3599
transform 1 0 15916 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_164
timestamp -3599
transform 1 0 16192 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_169
timestamp -3599
transform 1 0 16652 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_178
timestamp -3599
transform 1 0 17480 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_181
timestamp -3599
transform 1 0 17756 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_184
timestamp -3599
transform 1 0 18032 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_187
timestamp -3599
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_190
timestamp -3599
transform 1 0 18584 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_193
timestamp -3599
transform 1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_196
timestamp -3599
transform 1 0 19136 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_199
timestamp -3599
transform 1 0 19412 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_202
timestamp -3599
transform 1 0 19688 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_205
timestamp -3599
transform 1 0 19964 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_208
timestamp -3599
transform 1 0 20240 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_211
timestamp -3599
transform 1 0 20516 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_214
timestamp -3599
transform 1 0 20792 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_217
timestamp -3599
transform 1 0 21068 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_220
timestamp -3599
transform 1 0 21344 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp -3599
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp -3599
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_228
timestamp -3599
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_231
timestamp -3599
transform 1 0 22356 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_234
timestamp -3599
transform 1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_237
timestamp -3599
transform 1 0 22908 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_240
timestamp -3599
transform 1 0 23184 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_243
timestamp -3599
transform 1 0 23460 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_246
timestamp -3599
transform 1 0 23736 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_249
timestamp -3599
transform 1 0 24012 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_252
timestamp -3599
transform 1 0 24288 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_255
timestamp -3599
transform 1 0 24564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_258
timestamp -3599
transform 1 0 24840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_261
timestamp -3599
transform 1 0 25116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_264
timestamp -3599
transform 1 0 25392 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_267
timestamp -3599
transform 1 0 25668 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_270
timestamp -3599
transform 1 0 25944 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_273
timestamp -3599
transform 1 0 26220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_276
timestamp -3599
transform 1 0 26496 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp -3599
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_281
timestamp -3599
transform 1 0 26956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_284
timestamp -3599
transform 1 0 27232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_287
timestamp -3599
transform 1 0 27508 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_290
timestamp -3599
transform 1 0 27784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_293
timestamp -3599
transform 1 0 28060 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_296
timestamp -3599
transform 1 0 28336 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_299
timestamp -3599
transform 1 0 28612 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_303
timestamp -3599
transform 1 0 28980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_306
timestamp -3599
transform 1 0 29256 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_309
timestamp -3599
transform 1 0 29532 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_312
timestamp -3599
transform 1 0 29808 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_315
timestamp -3599
transform 1 0 30084 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_318
timestamp -3599
transform 1 0 30360 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_321
timestamp -3599
transform 1 0 30636 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_324
timestamp -3599
transform 1 0 30912 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_327
timestamp -3599
transform 1 0 31188 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_330
timestamp -3599
transform 1 0 31464 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_333
timestamp -3599
transform 1 0 31740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp -3599
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp -3599
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_6
timestamp -3599
transform 1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_9
timestamp -3599
transform 1 0 1932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_12
timestamp -3599
transform 1 0 2208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_15
timestamp -3599
transform 1 0 2484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_18
timestamp -3599
transform 1 0 2760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_21
timestamp -3599
transform 1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_24
timestamp -3599
transform 1 0 3312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -3599
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_29
timestamp -3599
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_32
timestamp -3599
transform 1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_35
timestamp -3599
transform 1 0 4324 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_38
timestamp -3599
transform 1 0 4600 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_41
timestamp -3599
transform 1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_44
timestamp -3599
transform 1 0 5152 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_47
timestamp -3599
transform 1 0 5428 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_50
timestamp -3599
transform 1 0 5704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_53
timestamp -3599
transform 1 0 5980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_56
timestamp -3599
transform 1 0 6256 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_59
timestamp -3599
transform 1 0 6532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_62
timestamp -3599
transform 1 0 6808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_65
timestamp -3599
transform 1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_68
timestamp -3599
transform 1 0 7360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_71
timestamp -3599
transform 1 0 7636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_74
timestamp -3599
transform 1 0 7912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_77
timestamp -3599
transform 1 0 8188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_80
timestamp -3599
transform 1 0 8464 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp -3599
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_85
timestamp -3599
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_88
timestamp -3599
transform 1 0 9200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_91
timestamp -3599
transform 1 0 9476 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_94
timestamp -3599
transform 1 0 9752 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_97
timestamp -3599
transform 1 0 10028 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_100
timestamp -3599
transform 1 0 10304 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_103
timestamp -3599
transform 1 0 10580 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_106
timestamp -3599
transform 1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_109
timestamp -3599
transform 1 0 11132 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_112
timestamp -3599
transform 1 0 11408 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_115
timestamp -3599
transform 1 0 11684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_118
timestamp -3599
transform 1 0 11960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_121
timestamp -3599
transform 1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_124
timestamp -3599
transform 1 0 12512 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_127
timestamp -3599
transform 1 0 12788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_130
timestamp -3599
transform 1 0 13064 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_133
timestamp -3599
transform 1 0 13340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_136
timestamp -3599
transform 1 0 13616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp -3599
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_141
timestamp -3599
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_144
timestamp -3599
transform 1 0 14352 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_147
timestamp -3599
transform 1 0 14628 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_150
timestamp -3599
transform 1 0 14904 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_153
timestamp -3599
transform 1 0 15180 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_156
timestamp -3599
transform 1 0 15456 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_159
timestamp -3599
transform 1 0 15732 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_162
timestamp -3599
transform 1 0 16008 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_165
timestamp -3599
transform 1 0 16284 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_168
timestamp -3599
transform 1 0 16560 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_171
timestamp -3599
transform 1 0 16836 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_183
timestamp -3599
transform 1 0 17940 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_186
timestamp -3599
transform 1 0 18216 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_189
timestamp -3599
transform 1 0 18492 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_192
timestamp -3599
transform 1 0 18768 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp -3599
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_197
timestamp -3599
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_200
timestamp -3599
transform 1 0 19504 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_203
timestamp -3599
transform 1 0 19780 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_206
timestamp -3599
transform 1 0 20056 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_209
timestamp -3599
transform 1 0 20332 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_212
timestamp -3599
transform 1 0 20608 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_215
timestamp -3599
transform 1 0 20884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_218
timestamp -3599
transform 1 0 21160 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_221
timestamp -3599
transform 1 0 21436 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_224
timestamp -3599
transform 1 0 21712 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_227
timestamp -3599
transform 1 0 21988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_230
timestamp -3599
transform 1 0 22264 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_233
timestamp -3599
transform 1 0 22540 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_236
timestamp -3599
transform 1 0 22816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_239
timestamp -3599
transform 1 0 23092 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_242
timestamp -3599
transform 1 0 23368 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_245
timestamp -3599
transform 1 0 23644 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_248
timestamp -3599
transform 1 0 23920 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp -3599
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp -3599
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_256
timestamp -3599
transform 1 0 24656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_259
timestamp -3599
transform 1 0 24932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_262
timestamp -3599
transform 1 0 25208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_265
timestamp -3599
transform 1 0 25484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_268
timestamp -3599
transform 1 0 25760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_271
timestamp -3599
transform 1 0 26036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_274
timestamp -3599
transform 1 0 26312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_277
timestamp -3599
transform 1 0 26588 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_280
timestamp -3599
transform 1 0 26864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_283
timestamp -3599
transform 1 0 27140 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_286
timestamp -3599
transform 1 0 27416 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_289
timestamp -3599
transform 1 0 27692 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_292
timestamp -3599
transform 1 0 27968 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_295
timestamp -3599
transform 1 0 28244 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_298
timestamp -3599
transform 1 0 28520 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_301
timestamp -3599
transform 1 0 28796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_304
timestamp -3599
transform 1 0 29072 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp -3599
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_309
timestamp -3599
transform 1 0 29532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_312
timestamp -3599
transform 1 0 29808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_315
timestamp -3599
transform 1 0 30084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_318
timestamp -3599
transform 1 0 30360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_321
timestamp -3599
transform 1 0 30636 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_326
timestamp -3599
transform 1 0 31096 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_329
timestamp -3599
transform 1 0 31372 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_332
timestamp -3599
transform 1 0 31648 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_335
timestamp -3599
transform 1 0 31924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_338
timestamp -3599
transform 1 0 32200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp -3599
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_6
timestamp -3599
transform 1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_9
timestamp -3599
transform 1 0 1932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_12
timestamp -3599
transform 1 0 2208 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_15
timestamp -3599
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_18
timestamp -3599
transform 1 0 2760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_21
timestamp -3599
transform 1 0 3036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_24
timestamp -3599
transform 1 0 3312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_27
timestamp -3599
transform 1 0 3588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_30
timestamp -3599
transform 1 0 3864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_33
timestamp -3599
transform 1 0 4140 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_36
timestamp -3599
transform 1 0 4416 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_39
timestamp -3599
transform 1 0 4692 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_42
timestamp -3599
transform 1 0 4968 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_45
timestamp -3599
transform 1 0 5244 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_48
timestamp -3599
transform 1 0 5520 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_51
timestamp -3599
transform 1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp -3599
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_57
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_60
timestamp -3599
transform 1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_63
timestamp -3599
transform 1 0 6900 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_66
timestamp -3599
transform 1 0 7176 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_69
timestamp -3599
transform 1 0 7452 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_72
timestamp -3599
transform 1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_75
timestamp -3599
transform 1 0 8004 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_78
timestamp -3599
transform 1 0 8280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_81
timestamp -3599
transform 1 0 8556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_84
timestamp -3599
transform 1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_87
timestamp -3599
transform 1 0 9108 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_90
timestamp -3599
transform 1 0 9384 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_93
timestamp -3599
transform 1 0 9660 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_96
timestamp -3599
transform 1 0 9936 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_99
timestamp -3599
transform 1 0 10212 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_102
timestamp -3599
transform 1 0 10488 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_105
timestamp -3599
transform 1 0 10764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_108
timestamp -3599
transform 1 0 11040 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp -3599
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_113
timestamp -3599
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_116
timestamp -3599
transform 1 0 11776 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_119
timestamp -3599
transform 1 0 12052 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_122
timestamp -3599
transform 1 0 12328 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_125
timestamp -3599
transform 1 0 12604 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_128
timestamp -3599
transform 1 0 12880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_131
timestamp -3599
transform 1 0 13156 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_134
timestamp -3599
transform 1 0 13432 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_137
timestamp -3599
transform 1 0 13708 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_140
timestamp -3599
transform 1 0 13984 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_143
timestamp -3599
transform 1 0 14260 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_146
timestamp -3599
transform 1 0 14536 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_149
timestamp -3599
transform 1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_152
timestamp -3599
transform 1 0 15088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_155
timestamp -3599
transform 1 0 15364 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_158
timestamp -3599
transform 1 0 15640 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_161
timestamp -3599
transform 1 0 15916 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_164
timestamp -3599
transform 1 0 16192 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp -3599
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_169
timestamp -3599
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_172
timestamp -3599
transform 1 0 16928 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_175
timestamp -3599
transform 1 0 17204 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_178
timestamp -3599
transform 1 0 17480 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_181
timestamp -3599
transform 1 0 17756 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_184
timestamp -3599
transform 1 0 18032 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_188
timestamp -3599
transform 1 0 18400 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_199
timestamp -3599
transform 1 0 19412 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_202
timestamp -3599
transform 1 0 19688 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_205
timestamp -3599
transform 1 0 19964 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_208
timestamp -3599
transform 1 0 20240 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_211
timestamp -3599
transform 1 0 20516 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_214
timestamp -3599
transform 1 0 20792 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_217
timestamp -3599
transform 1 0 21068 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_220
timestamp -3599
transform 1 0 21344 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp -3599
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp -3599
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_228
timestamp -3599
transform 1 0 22080 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_231
timestamp -3599
transform 1 0 22356 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_234
timestamp -3599
transform 1 0 22632 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_237
timestamp -3599
transform 1 0 22908 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_240
timestamp -3599
transform 1 0 23184 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_243
timestamp -3599
transform 1 0 23460 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_246
timestamp -3599
transform 1 0 23736 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_249
timestamp -3599
transform 1 0 24012 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_252
timestamp -3599
transform 1 0 24288 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_255
timestamp -3599
transform 1 0 24564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_258
timestamp -3599
transform 1 0 24840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_261
timestamp -3599
transform 1 0 25116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_264
timestamp -3599
transform 1 0 25392 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_267
timestamp -3599
transform 1 0 25668 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_270
timestamp -3599
transform 1 0 25944 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_273
timestamp -3599
transform 1 0 26220 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_276
timestamp -3599
transform 1 0 26496 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp -3599
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_281
timestamp -3599
transform 1 0 26956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_284
timestamp -3599
transform 1 0 27232 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_287
timestamp -3599
transform 1 0 27508 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_290
timestamp -3599
transform 1 0 27784 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_293
timestamp -3599
transform 1 0 28060 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_296
timestamp -3599
transform 1 0 28336 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_299
timestamp -3599
transform 1 0 28612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_302
timestamp -3599
transform 1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_305
timestamp -3599
transform 1 0 29164 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_308
timestamp -3599
transform 1 0 29440 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_314
timestamp -3599
transform 1 0 29992 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_317
timestamp -3599
transform 1 0 30268 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_320
timestamp -3599
transform 1 0 30544 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_323
timestamp -3599
transform 1 0 30820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_326
timestamp -3599
transform 1 0 31096 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_329
timestamp -3599
transform 1 0 31372 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_332
timestamp -3599
transform 1 0 31648 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp -3599
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp -3599
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_6
timestamp -3599
transform 1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_9
timestamp -3599
transform 1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_12
timestamp -3599
transform 1 0 2208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_15
timestamp -3599
transform 1 0 2484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_18
timestamp -3599
transform 1 0 2760 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_21
timestamp -3599
transform 1 0 3036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_24
timestamp -3599
transform 1 0 3312 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp -3599
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_29
timestamp -3599
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_32
timestamp -3599
transform 1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_35
timestamp -3599
transform 1 0 4324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_38
timestamp -3599
transform 1 0 4600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_41
timestamp -3599
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_44
timestamp -3599
transform 1 0 5152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_47
timestamp -3599
transform 1 0 5428 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_50
timestamp -3599
transform 1 0 5704 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_53
timestamp -3599
transform 1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_56
timestamp -3599
transform 1 0 6256 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_59
timestamp -3599
transform 1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_62
timestamp -3599
transform 1 0 6808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_65
timestamp -3599
transform 1 0 7084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_68
timestamp -3599
transform 1 0 7360 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_71
timestamp -3599
transform 1 0 7636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_74
timestamp -3599
transform 1 0 7912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_77
timestamp -3599
transform 1 0 8188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_80
timestamp -3599
transform 1 0 8464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp -3599
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_85
timestamp -3599
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_88
timestamp -3599
transform 1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_91
timestamp -3599
transform 1 0 9476 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_94
timestamp -3599
transform 1 0 9752 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_97
timestamp -3599
transform 1 0 10028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_100
timestamp -3599
transform 1 0 10304 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_103
timestamp -3599
transform 1 0 10580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_106
timestamp -3599
transform 1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_109
timestamp -3599
transform 1 0 11132 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_112
timestamp -3599
transform 1 0 11408 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_115
timestamp -3599
transform 1 0 11684 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_118
timestamp -3599
transform 1 0 11960 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_121
timestamp -3599
transform 1 0 12236 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_124
timestamp -3599
transform 1 0 12512 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_127
timestamp -3599
transform 1 0 12788 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_130
timestamp -3599
transform 1 0 13064 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_133
timestamp -3599
transform 1 0 13340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_136
timestamp -3599
transform 1 0 13616 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp -3599
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_141
timestamp -3599
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_144
timestamp -3599
transform 1 0 14352 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_147
timestamp -3599
transform 1 0 14628 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_150
timestamp -3599
transform 1 0 14904 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_153
timestamp -3599
transform 1 0 15180 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_156
timestamp -3599
transform 1 0 15456 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_159
timestamp -3599
transform 1 0 15732 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_162
timestamp -3599
transform 1 0 16008 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_165
timestamp -3599
transform 1 0 16284 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_168
timestamp -3599
transform 1 0 16560 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_171
timestamp -3599
transform 1 0 16836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_174
timestamp -3599
transform 1 0 17112 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_177
timestamp -3599
transform 1 0 17388 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_180
timestamp -3599
transform 1 0 17664 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_183
timestamp -3599
transform 1 0 17940 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_186
timestamp -3599
transform 1 0 18216 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_189
timestamp -3599
transform 1 0 18492 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_192
timestamp -3599
transform 1 0 18768 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp -3599
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp -3599
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_200
timestamp -3599
transform 1 0 19504 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_203
timestamp -3599
transform 1 0 19780 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_206
timestamp -3599
transform 1 0 20056 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_211
timestamp -3599
transform 1 0 20516 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_215
timestamp -3599
transform 1 0 20884 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_224
timestamp -3599
transform 1 0 21712 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_227
timestamp -3599
transform 1 0 21988 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_230
timestamp -3599
transform 1 0 22264 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_233
timestamp -3599
transform 1 0 22540 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_236
timestamp -3599
transform 1 0 22816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_239
timestamp -3599
transform 1 0 23092 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_242
timestamp -3599
transform 1 0 23368 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_245
timestamp -3599
transform 1 0 23644 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_248
timestamp -3599
transform 1 0 23920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp -3599
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_259
timestamp -3599
transform 1 0 24932 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_264
timestamp -3599
transform 1 0 25392 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_267
timestamp -3599
transform 1 0 25668 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_270
timestamp -3599
transform 1 0 25944 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_274
timestamp -3599
transform 1 0 26312 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_277
timestamp -3599
transform 1 0 26588 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_280
timestamp -3599
transform 1 0 26864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_283
timestamp -3599
transform 1 0 27140 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_286
timestamp -3599
transform 1 0 27416 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_289
timestamp -3599
transform 1 0 27692 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_292
timestamp -3599
transform 1 0 27968 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_295
timestamp -3599
transform 1 0 28244 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_298
timestamp -3599
transform 1 0 28520 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_303
timestamp -3599
transform 1 0 28980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp -3599
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_309
timestamp -3599
transform 1 0 29532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_312
timestamp -3599
transform 1 0 29808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_315
timestamp -3599
transform 1 0 30084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_318
timestamp -3599
transform 1 0 30360 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_321
timestamp -3599
transform 1 0 30636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_324
timestamp -3599
transform 1 0 30912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_327
timestamp -3599
transform 1 0 31188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_330
timestamp -3599
transform 1 0 31464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_333
timestamp -3599
transform 1 0 31740 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_336
timestamp -3599
transform 1 0 32016 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp -3599
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6
timestamp -3599
transform 1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_9
timestamp -3599
transform 1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_12
timestamp -3599
transform 1 0 2208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_15
timestamp -3599
transform 1 0 2484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_18
timestamp -3599
transform 1 0 2760 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_21
timestamp -3599
transform 1 0 3036 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_24
timestamp -3599
transform 1 0 3312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_27
timestamp -3599
transform 1 0 3588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_30
timestamp -3599
transform 1 0 3864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_33
timestamp -3599
transform 1 0 4140 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_36
timestamp -3599
transform 1 0 4416 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_39
timestamp -3599
transform 1 0 4692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_42
timestamp -3599
transform 1 0 4968 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_45
timestamp -3599
transform 1 0 5244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_48
timestamp -3599
transform 1 0 5520 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_51
timestamp -3599
transform 1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp -3599
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp -3599
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_60
timestamp -3599
transform 1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_63
timestamp -3599
transform 1 0 6900 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_66
timestamp -3599
transform 1 0 7176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_69
timestamp -3599
transform 1 0 7452 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_72
timestamp -3599
transform 1 0 7728 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_75
timestamp -3599
transform 1 0 8004 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_78
timestamp -3599
transform 1 0 8280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_81
timestamp -3599
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_84
timestamp -3599
transform 1 0 8832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_92
timestamp -3599
transform 1 0 9568 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_95
timestamp -3599
transform 1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_98
timestamp -3599
transform 1 0 10120 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_101
timestamp -3599
transform 1 0 10396 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_104
timestamp -3599
transform 1 0 10672 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp -3599
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_113
timestamp -3599
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_116
timestamp -3599
transform 1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_119
timestamp -3599
transform 1 0 12052 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_123
timestamp -3599
transform 1 0 12420 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_126
timestamp -3599
transform 1 0 12696 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_129
timestamp -3599
transform 1 0 12972 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_132
timestamp -3599
transform 1 0 13248 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_135
timestamp -3599
transform 1 0 13524 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_138
timestamp -3599
transform 1 0 13800 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_141
timestamp -3599
transform 1 0 14076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_145
timestamp -3599
transform 1 0 14444 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_152
timestamp -3599
transform 1 0 15088 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_155
timestamp -3599
transform 1 0 15364 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_158
timestamp -3599
transform 1 0 15640 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_161
timestamp -3599
transform 1 0 15916 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_164
timestamp -3599
transform 1 0 16192 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp -3599
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_169
timestamp -3599
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_172
timestamp -3599
transform 1 0 16928 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_175
timestamp -3599
transform 1 0 17204 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_178
timestamp -3599
transform 1 0 17480 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_187
timestamp -3599
transform 1 0 18308 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_190
timestamp -3599
transform 1 0 18584 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_193
timestamp -3599
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_196
timestamp -3599
transform 1 0 19136 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_199
timestamp -3599
transform 1 0 19412 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_202
timestamp -3599
transform 1 0 19688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_206
timestamp -3599
transform 1 0 20056 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_209
timestamp -3599
transform 1 0 20332 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_212
timestamp -3599
transform 1 0 20608 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_215
timestamp -3599
transform 1 0 20884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_218
timestamp -3599
transform 1 0 21160 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp -3599
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_228
timestamp -3599
transform 1 0 22080 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_235
timestamp -3599
transform 1 0 22724 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_238
timestamp -3599
transform 1 0 23000 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_241
timestamp -3599
transform 1 0 23276 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_244
timestamp -3599
transform 1 0 23552 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_247
timestamp -3599
transform 1 0 23828 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_260
timestamp -3599
transform 1 0 25024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_266
timestamp -3599
transform 1 0 25576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_269
timestamp -3599
transform 1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_272
timestamp -3599
transform 1 0 26128 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_275
timestamp -3599
transform 1 0 26404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp -3599
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_281
timestamp -3599
transform 1 0 26956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_284
timestamp -3599
transform 1 0 27232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_287
timestamp -3599
transform 1 0 27508 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_301
timestamp -3599
transform 1 0 28796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_304
timestamp -3599
transform 1 0 29072 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_307
timestamp -3599
transform 1 0 29348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_311
timestamp -3599
transform 1 0 29716 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_314
timestamp -3599
transform 1 0 29992 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_317
timestamp -3599
transform 1 0 30268 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_320
timestamp -3599
transform 1 0 30544 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_323
timestamp -3599
transform 1 0 30820 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_327
timestamp -3599
transform 1 0 31188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_330
timestamp -3599
transform 1 0 31464 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp -3599
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp -3599
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_6
timestamp -3599
transform 1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_9
timestamp -3599
transform 1 0 1932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_12
timestamp -3599
transform 1 0 2208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_15
timestamp -3599
transform 1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_18
timestamp -3599
transform 1 0 2760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_21
timestamp -3599
transform 1 0 3036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_24
timestamp -3599
transform 1 0 3312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp -3599
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_32
timestamp -3599
transform 1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_35
timestamp -3599
transform 1 0 4324 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_38
timestamp -3599
transform 1 0 4600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_41
timestamp -3599
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_44
timestamp -3599
transform 1 0 5152 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_47
timestamp -3599
transform 1 0 5428 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_50
timestamp -3599
transform 1 0 5704 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_53
timestamp -3599
transform 1 0 5980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_56
timestamp -3599
transform 1 0 6256 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_59
timestamp -3599
transform 1 0 6532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_62
timestamp -3599
transform 1 0 6808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_65
timestamp -3599
transform 1 0 7084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_68
timestamp -3599
transform 1 0 7360 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_71
timestamp -3599
transform 1 0 7636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_74
timestamp -3599
transform 1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_77
timestamp -3599
transform 1 0 8188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_80
timestamp -3599
transform 1 0 8464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp -3599
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_85
timestamp -3599
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_88
timestamp -3599
transform 1 0 9200 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_91
timestamp -3599
transform 1 0 9476 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_94
timestamp -3599
transform 1 0 9752 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_97
timestamp -3599
transform 1 0 10028 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_100
timestamp -3599
transform 1 0 10304 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_103
timestamp -3599
transform 1 0 10580 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_106
timestamp -3599
transform 1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_109
timestamp -3599
transform 1 0 11132 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_112
timestamp -3599
transform 1 0 11408 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_115
timestamp -3599
transform 1 0 11684 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_118
timestamp -3599
transform 1 0 11960 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_121
timestamp -3599
transform 1 0 12236 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_124
timestamp -3599
transform 1 0 12512 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_127
timestamp -3599
transform 1 0 12788 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_130
timestamp -3599
transform 1 0 13064 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_133
timestamp -3599
transform 1 0 13340 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_136
timestamp -3599
transform 1 0 13616 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp -3599
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_141
timestamp -3599
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_144
timestamp -3599
transform 1 0 14352 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_147
timestamp -3599
transform 1 0 14628 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_150
timestamp -3599
transform 1 0 14904 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_153
timestamp -3599
transform 1 0 15180 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_156
timestamp -3599
transform 1 0 15456 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_159
timestamp -3599
transform 1 0 15732 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_162
timestamp -3599
transform 1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_165
timestamp -3599
transform 1 0 16284 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_168
timestamp -3599
transform 1 0 16560 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_171
timestamp -3599
transform 1 0 16836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_174
timestamp -3599
transform 1 0 17112 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_177
timestamp -3599
transform 1 0 17388 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_180
timestamp -3599
transform 1 0 17664 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_183
timestamp -3599
transform 1 0 17940 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_186
timestamp -3599
transform 1 0 18216 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_189
timestamp -3599
transform 1 0 18492 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_192
timestamp -3599
transform 1 0 18768 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp -3599
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_197
timestamp -3599
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_200
timestamp -3599
transform 1 0 19504 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_203
timestamp -3599
transform 1 0 19780 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_206
timestamp -3599
transform 1 0 20056 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_209
timestamp -3599
transform 1 0 20332 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_212
timestamp -3599
transform 1 0 20608 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_215
timestamp -3599
transform 1 0 20884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_218
timestamp -3599
transform 1 0 21160 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_221
timestamp -3599
transform 1 0 21436 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_224
timestamp -3599
transform 1 0 21712 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_227
timestamp -3599
transform 1 0 21988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_230
timestamp -3599
transform 1 0 22264 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_233
timestamp -3599
transform 1 0 22540 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_236
timestamp -3599
transform 1 0 22816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_239
timestamp -3599
transform 1 0 23092 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_242
timestamp -3599
transform 1 0 23368 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_245
timestamp -3599
transform 1 0 23644 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_248
timestamp -3599
transform 1 0 23920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp -3599
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_253
timestamp -3599
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_256
timestamp -3599
transform 1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_259
timestamp -3599
transform 1 0 24932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_262
timestamp -3599
transform 1 0 25208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_265
timestamp -3599
transform 1 0 25484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_268
timestamp -3599
transform 1 0 25760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_271
timestamp -3599
transform 1 0 26036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_274
timestamp -3599
transform 1 0 26312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_277
timestamp -3599
transform 1 0 26588 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_280
timestamp -3599
transform 1 0 26864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_283
timestamp -3599
transform 1 0 27140 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_286
timestamp -3599
transform 1 0 27416 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_289
timestamp -3599
transform 1 0 27692 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_292
timestamp -3599
transform 1 0 27968 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_295
timestamp -3599
transform 1 0 28244 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_298
timestamp -3599
transform 1 0 28520 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_301
timestamp -3599
transform 1 0 28796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_304
timestamp -3599
transform 1 0 29072 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp -3599
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_309
timestamp -3599
transform 1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_312
timestamp -3599
transform 1 0 29808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_315
timestamp -3599
transform 1 0 30084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_318
timestamp -3599
transform 1 0 30360 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_321
timestamp -3599
transform 1 0 30636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_324
timestamp -3599
transform 1 0 30912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp -3599
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_8
timestamp -3599
transform 1 0 1840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_11
timestamp -3599
transform 1 0 2116 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_14
timestamp -3599
transform 1 0 2392 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_17
timestamp -3599
transform 1 0 2668 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_20
timestamp -3599
transform 1 0 2944 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_26
timestamp -3599
transform 1 0 3496 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_29
timestamp -3599
transform 1 0 3772 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_32
timestamp -3599
transform 1 0 4048 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_35
timestamp -3599
transform 1 0 4324 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_38
timestamp -3599
transform 1 0 4600 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_43
timestamp -3599
transform 1 0 5060 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_46
timestamp -3599
transform 1 0 5336 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_49
timestamp -3599
transform 1 0 5612 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_52
timestamp -3599
transform 1 0 5888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp -3599
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_61
timestamp -3599
transform 1 0 6716 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_64
timestamp -3599
transform 1 0 6992 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_67
timestamp -3599
transform 1 0 7268 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_70
timestamp -3599
transform 1 0 7544 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_77
timestamp -3599
transform 1 0 8188 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_80
timestamp -3599
transform 1 0 8464 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_83
timestamp -3599
transform 1 0 8740 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_85
timestamp -3599
transform 1 0 8924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_88
timestamp -3599
transform 1 0 9200 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_94
timestamp -3599
transform 1 0 9752 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_97
timestamp -3599
transform 1 0 10028 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_100
timestamp -3599
transform 1 0 10304 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_103
timestamp -3599
transform 1 0 10580 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_106
timestamp -3599
transform 1 0 10856 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp -3599
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp -3599
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_116
timestamp -3599
transform 1 0 11776 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_119
timestamp -3599
transform 1 0 12052 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_122
timestamp -3599
transform 1 0 12328 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_128
timestamp -3599
transform 1 0 12880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_131
timestamp -3599
transform 1 0 13156 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_134
timestamp -3599
transform 1 0 13432 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_137
timestamp -3599
transform 1 0 13708 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_145
timestamp -3599
transform 1 0 14444 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_148
timestamp -3599
transform 1 0 14720 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_151
timestamp -3599
transform 1 0 14996 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_154
timestamp -3599
transform 1 0 15272 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_157
timestamp -3599
transform 1 0 15548 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_162
timestamp -3599
transform 1 0 16008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp -3599
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp -3599
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_172
timestamp -3599
transform 1 0 16928 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_179
timestamp -3599
transform 1 0 17572 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_182
timestamp -3599
transform 1 0 17848 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_185
timestamp -3599
transform 1 0 18124 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_188
timestamp -3599
transform 1 0 18400 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_191
timestamp -3599
transform 1 0 18676 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_197
timestamp -3599
transform 1 0 19228 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_200
timestamp -3599
transform 1 0 19504 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_203
timestamp -3599
transform 1 0 19780 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_206
timestamp -3599
transform 1 0 20056 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_213
timestamp -3599
transform 1 0 20700 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_216
timestamp -3599
transform 1 0 20976 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_219
timestamp -3599
transform 1 0 21252 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp -3599
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_225
timestamp -3599
transform 1 0 21804 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_230
timestamp -3599
transform 1 0 22264 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_233
timestamp -3599
transform 1 0 22540 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_236
timestamp -3599
transform 1 0 22816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_239
timestamp -3599
transform 1 0 23092 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_242
timestamp -3599
transform 1 0 23368 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_247
timestamp -3599
transform 1 0 23828 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_250
timestamp -3599
transform 1 0 24104 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_253
timestamp -3599
transform 1 0 24380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_256
timestamp -3599
transform 1 0 24656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_259
timestamp -3599
transform 1 0 24932 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_264
timestamp -3599
transform 1 0 25392 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_267
timestamp -3599
transform 1 0 25668 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_270
timestamp -3599
transform 1 0 25944 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_273
timestamp -3599
transform 1 0 26220 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_276
timestamp -3599
transform 1 0 26496 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp -3599
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_285
timestamp -3599
transform 1 0 27324 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_288
timestamp -3599
transform 1 0 27600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_291
timestamp -3599
transform 1 0 27876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_298
timestamp -3599
transform 1 0 28520 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_301
timestamp -3599
transform 1 0 28796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_304
timestamp -3599
transform 1 0 29072 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_307
timestamp -3599
transform 1 0 29348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_309
timestamp -3599
transform 1 0 29532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_315
timestamp -3599
transform 1 0 30084 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_318
timestamp -3599
transform 1 0 30360 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_321
timestamp -3599
transform 1 0 30636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp -3599
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output1
timestamp -3599
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp -3599
transform 1 0 32292 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp -3599
transform 1 0 32660 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp -3599
transform 1 0 32292 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp -3599
transform 1 0 32660 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp -3599
transform 1 0 32292 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp -3599
transform 1 0 32660 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp -3599
transform 1 0 32292 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp -3599
transform 1 0 32660 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp -3599
transform 1 0 32292 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp -3599
transform 1 0 32660 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp -3599
transform 1 0 31280 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp -3599
transform 1 0 32292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp -3599
transform 1 0 32660 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp -3599
transform 1 0 32660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp -3599
transform 1 0 32292 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp -3599
transform 1 0 32660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp -3599
transform 1 0 32292 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp -3599
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp -3599
transform 1 0 31924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp -3599
transform 1 0 32292 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp -3599
transform 1 0 31556 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp -3599
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp -3599
transform 1 0 30912 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp -3599
transform 1 0 31188 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp -3599
transform 1 0 30912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp -3599
transform 1 0 32292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp -3599
transform 1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp -3599
transform 1 0 32292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp -3599
transform 1 0 32660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp -3599
transform 1 0 32292 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp -3599
transform 1 0 32660 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp -3599
transform -1 0 3496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp -3599
transform -1 0 19136 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp -3599
transform -1 0 20700 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp -3599
transform -1 0 22264 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp -3599
transform -1 0 23828 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp -3599
transform 1 0 25024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp -3599
transform -1 0 27324 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp -3599
transform -1 0 28520 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp -3599
transform 1 0 29716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp -3599
transform 1 0 31280 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp -3599
transform 1 0 32660 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp -3599
transform -1 0 5060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp -3599
transform -1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp -3599
transform -1 0 8188 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp -3599
transform -1 0 9752 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp -3599
transform -1 0 11316 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp -3599
transform -1 0 12880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp -3599
transform -1 0 14444 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp -3599
transform -1 0 16008 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp -3599
transform -1 0 17572 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp -3599
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp -3599
transform 1 0 14720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp -3599
transform 1 0 15824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp -3599
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp -3599
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp -3599
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp -3599
transform 1 0 15824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp -3599
transform 1 0 16744 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp -3599
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp -3599
transform 1 0 17112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp -3599
transform 1 0 16928 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp -3599
transform 1 0 17480 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp -3599
transform 1 0 17296 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp -3599
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp -3599
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp -3599
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp -3599
transform 1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp -3599
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp -3599
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp -3599
transform 1 0 18952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp -3599
transform 1 0 19964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp -3599
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp -3599
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp -3599
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp -3599
transform 1 0 22540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp -3599
transform 1 0 22172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp -3599
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp -3599
transform 1 0 19320 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp -3599
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp -3599
transform 1 0 19688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp -3599
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp -3599
transform 1 0 20056 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp -3599
transform 1 0 21068 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp -3599
transform 1 0 20424 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp -3599
transform 1 0 20792 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform 1 0 21160 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp -3599
transform -1 0 22908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp -3599
transform -1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp -3599
transform -1 0 25116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp -3599
transform -1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp -3599
transform -1 0 25484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp -3599
transform -1 0 26220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp -3599
transform -1 0 25852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp -3599
transform -1 0 23644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp -3599
transform -1 0 23276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp -3599
transform -1 0 24012 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp -3599
transform -1 0 23644 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp -3599
transform -1 0 24012 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp -3599
transform -1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp -3599
transform -1 0 24380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp -3599
transform -1 0 25116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp -3599
transform -1 0 24748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output105
timestamp -3599
transform -1 0 1840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 33304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 33304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 33304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 33304 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 33304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 33304 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 33304 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 33304 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 33304 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 33304 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 33304 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 33304 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp -3599
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp -3599
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_36
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_37
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_38
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_39
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_40
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_41
timestamp -3599
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_42
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_43
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_44
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_45
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_46
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_47
timestamp -3599
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_48
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_49
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_50
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_51
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_52
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_53
timestamp -3599
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_54
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_55
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_56
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_57
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_58
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_59
timestamp -3599
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_60
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_61
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_62
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_63
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_64
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_65
timestamp -3599
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_66
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_67
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_68
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_69
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_70
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_71
timestamp -3599
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_72
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_73
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_74
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_75
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_76
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_77
timestamp -3599
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_78
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_79
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_80
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_81
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_82
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_83
timestamp -3599
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_84
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_85
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_86
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_87
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_88
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_89
timestamp -3599
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_90
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_91
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_92
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_93
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_94
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_95
timestamp -3599
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_96
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_97
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_98
timestamp -3599
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_99
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_100
timestamp -3599
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_101
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_102
timestamp -3599
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_103
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_104
timestamp -3599
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_105
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_106
timestamp -3599
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_107
timestamp -3599
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 15198 0 15254 56 0 FreeSans 224 0 0 0 Ci
port 0 nsew signal input
flabel metal3 s 0 1096 120 1216 0 FreeSans 480 0 0 0 FrameData[0]
port 1 nsew signal input
flabel metal3 s 0 3816 120 3936 0 FreeSans 480 0 0 0 FrameData[10]
port 2 nsew signal input
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 FrameData[11]
port 3 nsew signal input
flabel metal3 s 0 4360 120 4480 0 FreeSans 480 0 0 0 FrameData[12]
port 4 nsew signal input
flabel metal3 s 0 4632 120 4752 0 FreeSans 480 0 0 0 FrameData[13]
port 5 nsew signal input
flabel metal3 s 0 4904 120 5024 0 FreeSans 480 0 0 0 FrameData[14]
port 6 nsew signal input
flabel metal3 s 0 5176 120 5296 0 FreeSans 480 0 0 0 FrameData[15]
port 7 nsew signal input
flabel metal3 s 0 5448 120 5568 0 FreeSans 480 0 0 0 FrameData[16]
port 8 nsew signal input
flabel metal3 s 0 5720 120 5840 0 FreeSans 480 0 0 0 FrameData[17]
port 9 nsew signal input
flabel metal3 s 0 5992 120 6112 0 FreeSans 480 0 0 0 FrameData[18]
port 10 nsew signal input
flabel metal3 s 0 6264 120 6384 0 FreeSans 480 0 0 0 FrameData[19]
port 11 nsew signal input
flabel metal3 s 0 1368 120 1488 0 FreeSans 480 0 0 0 FrameData[1]
port 12 nsew signal input
flabel metal3 s 0 6536 120 6656 0 FreeSans 480 0 0 0 FrameData[20]
port 13 nsew signal input
flabel metal3 s 0 6808 120 6928 0 FreeSans 480 0 0 0 FrameData[21]
port 14 nsew signal input
flabel metal3 s 0 7080 120 7200 0 FreeSans 480 0 0 0 FrameData[22]
port 15 nsew signal input
flabel metal3 s 0 7352 120 7472 0 FreeSans 480 0 0 0 FrameData[23]
port 16 nsew signal input
flabel metal3 s 0 7624 120 7744 0 FreeSans 480 0 0 0 FrameData[24]
port 17 nsew signal input
flabel metal3 s 0 7896 120 8016 0 FreeSans 480 0 0 0 FrameData[25]
port 18 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 FrameData[26]
port 19 nsew signal input
flabel metal3 s 0 8440 120 8560 0 FreeSans 480 0 0 0 FrameData[27]
port 20 nsew signal input
flabel metal3 s 0 8712 120 8832 0 FreeSans 480 0 0 0 FrameData[28]
port 21 nsew signal input
flabel metal3 s 0 8984 120 9104 0 FreeSans 480 0 0 0 FrameData[29]
port 22 nsew signal input
flabel metal3 s 0 1640 120 1760 0 FreeSans 480 0 0 0 FrameData[2]
port 23 nsew signal input
flabel metal3 s 0 9256 120 9376 0 FreeSans 480 0 0 0 FrameData[30]
port 24 nsew signal input
flabel metal3 s 0 9528 120 9648 0 FreeSans 480 0 0 0 FrameData[31]
port 25 nsew signal input
flabel metal3 s 0 1912 120 2032 0 FreeSans 480 0 0 0 FrameData[3]
port 26 nsew signal input
flabel metal3 s 0 2184 120 2304 0 FreeSans 480 0 0 0 FrameData[4]
port 27 nsew signal input
flabel metal3 s 0 2456 120 2576 0 FreeSans 480 0 0 0 FrameData[5]
port 28 nsew signal input
flabel metal3 s 0 2728 120 2848 0 FreeSans 480 0 0 0 FrameData[6]
port 29 nsew signal input
flabel metal3 s 0 3000 120 3120 0 FreeSans 480 0 0 0 FrameData[7]
port 30 nsew signal input
flabel metal3 s 0 3272 120 3392 0 FreeSans 480 0 0 0 FrameData[8]
port 31 nsew signal input
flabel metal3 s 0 3544 120 3664 0 FreeSans 480 0 0 0 FrameData[9]
port 32 nsew signal input
flabel metal3 s 34288 1096 34408 1216 0 FreeSans 480 0 0 0 FrameData_O[0]
port 33 nsew signal output
flabel metal3 s 34288 3816 34408 3936 0 FreeSans 480 0 0 0 FrameData_O[10]
port 34 nsew signal output
flabel metal3 s 34288 4088 34408 4208 0 FreeSans 480 0 0 0 FrameData_O[11]
port 35 nsew signal output
flabel metal3 s 34288 4360 34408 4480 0 FreeSans 480 0 0 0 FrameData_O[12]
port 36 nsew signal output
flabel metal3 s 34288 4632 34408 4752 0 FreeSans 480 0 0 0 FrameData_O[13]
port 37 nsew signal output
flabel metal3 s 34288 4904 34408 5024 0 FreeSans 480 0 0 0 FrameData_O[14]
port 38 nsew signal output
flabel metal3 s 34288 5176 34408 5296 0 FreeSans 480 0 0 0 FrameData_O[15]
port 39 nsew signal output
flabel metal3 s 34288 5448 34408 5568 0 FreeSans 480 0 0 0 FrameData_O[16]
port 40 nsew signal output
flabel metal3 s 34288 5720 34408 5840 0 FreeSans 480 0 0 0 FrameData_O[17]
port 41 nsew signal output
flabel metal3 s 34288 5992 34408 6112 0 FreeSans 480 0 0 0 FrameData_O[18]
port 42 nsew signal output
flabel metal3 s 34288 6264 34408 6384 0 FreeSans 480 0 0 0 FrameData_O[19]
port 43 nsew signal output
flabel metal3 s 34288 1368 34408 1488 0 FreeSans 480 0 0 0 FrameData_O[1]
port 44 nsew signal output
flabel metal3 s 34288 6536 34408 6656 0 FreeSans 480 0 0 0 FrameData_O[20]
port 45 nsew signal output
flabel metal3 s 34288 6808 34408 6928 0 FreeSans 480 0 0 0 FrameData_O[21]
port 46 nsew signal output
flabel metal3 s 34288 7080 34408 7200 0 FreeSans 480 0 0 0 FrameData_O[22]
port 47 nsew signal output
flabel metal3 s 34288 7352 34408 7472 0 FreeSans 480 0 0 0 FrameData_O[23]
port 48 nsew signal output
flabel metal3 s 34288 7624 34408 7744 0 FreeSans 480 0 0 0 FrameData_O[24]
port 49 nsew signal output
flabel metal3 s 34288 7896 34408 8016 0 FreeSans 480 0 0 0 FrameData_O[25]
port 50 nsew signal output
flabel metal3 s 34288 8168 34408 8288 0 FreeSans 480 0 0 0 FrameData_O[26]
port 51 nsew signal output
flabel metal3 s 34288 8440 34408 8560 0 FreeSans 480 0 0 0 FrameData_O[27]
port 52 nsew signal output
flabel metal3 s 34288 8712 34408 8832 0 FreeSans 480 0 0 0 FrameData_O[28]
port 53 nsew signal output
flabel metal3 s 34288 8984 34408 9104 0 FreeSans 480 0 0 0 FrameData_O[29]
port 54 nsew signal output
flabel metal3 s 34288 1640 34408 1760 0 FreeSans 480 0 0 0 FrameData_O[2]
port 55 nsew signal output
flabel metal3 s 34288 9256 34408 9376 0 FreeSans 480 0 0 0 FrameData_O[30]
port 56 nsew signal output
flabel metal3 s 34288 9528 34408 9648 0 FreeSans 480 0 0 0 FrameData_O[31]
port 57 nsew signal output
flabel metal3 s 34288 1912 34408 2032 0 FreeSans 480 0 0 0 FrameData_O[3]
port 58 nsew signal output
flabel metal3 s 34288 2184 34408 2304 0 FreeSans 480 0 0 0 FrameData_O[4]
port 59 nsew signal output
flabel metal3 s 34288 2456 34408 2576 0 FreeSans 480 0 0 0 FrameData_O[5]
port 60 nsew signal output
flabel metal3 s 34288 2728 34408 2848 0 FreeSans 480 0 0 0 FrameData_O[6]
port 61 nsew signal output
flabel metal3 s 34288 3000 34408 3120 0 FreeSans 480 0 0 0 FrameData_O[7]
port 62 nsew signal output
flabel metal3 s 34288 3272 34408 3392 0 FreeSans 480 0 0 0 FrameData_O[8]
port 63 nsew signal output
flabel metal3 s 34288 3544 34408 3664 0 FreeSans 480 0 0 0 FrameData_O[9]
port 64 nsew signal output
flabel metal2 s 25134 0 25190 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 65 nsew signal input
flabel metal2 s 26974 0 27030 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 66 nsew signal input
flabel metal2 s 27158 0 27214 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 67 nsew signal input
flabel metal2 s 27342 0 27398 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 68 nsew signal input
flabel metal2 s 27526 0 27582 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 69 nsew signal input
flabel metal2 s 27710 0 27766 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 70 nsew signal input
flabel metal2 s 27894 0 27950 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 71 nsew signal input
flabel metal2 s 28078 0 28134 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 72 nsew signal input
flabel metal2 s 28262 0 28318 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 73 nsew signal input
flabel metal2 s 28446 0 28502 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 74 nsew signal input
flabel metal2 s 28630 0 28686 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 75 nsew signal input
flabel metal2 s 25318 0 25374 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 76 nsew signal input
flabel metal2 s 25502 0 25558 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 77 nsew signal input
flabel metal2 s 25686 0 25742 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 78 nsew signal input
flabel metal2 s 25870 0 25926 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 79 nsew signal input
flabel metal2 s 26054 0 26110 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 80 nsew signal input
flabel metal2 s 26238 0 26294 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 81 nsew signal input
flabel metal2 s 26422 0 26478 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 82 nsew signal input
flabel metal2 s 26606 0 26662 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 83 nsew signal input
flabel metal2 s 26790 0 26846 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 84 nsew signal input
flabel metal2 s 3054 11096 3110 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 85 nsew signal output
flabel metal2 s 18694 11096 18750 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 86 nsew signal output
flabel metal2 s 20258 11096 20314 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 87 nsew signal output
flabel metal2 s 21822 11096 21878 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 88 nsew signal output
flabel metal2 s 23386 11096 23442 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 89 nsew signal output
flabel metal2 s 24950 11096 25006 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 90 nsew signal output
flabel metal2 s 26514 11096 26570 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 91 nsew signal output
flabel metal2 s 28078 11096 28134 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 92 nsew signal output
flabel metal2 s 29642 11096 29698 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 93 nsew signal output
flabel metal2 s 31206 11096 31262 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 94 nsew signal output
flabel metal2 s 32770 11096 32826 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 95 nsew signal output
flabel metal2 s 4618 11096 4674 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 96 nsew signal output
flabel metal2 s 6182 11096 6238 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 97 nsew signal output
flabel metal2 s 7746 11096 7802 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 98 nsew signal output
flabel metal2 s 9310 11096 9366 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 99 nsew signal output
flabel metal2 s 10874 11096 10930 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 100 nsew signal output
flabel metal2 s 12438 11096 12494 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 101 nsew signal output
flabel metal2 s 14002 11096 14058 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 102 nsew signal output
flabel metal2 s 15566 11096 15622 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 103 nsew signal output
flabel metal2 s 17130 11096 17186 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 104 nsew signal output
flabel metal2 s 5630 0 5686 56 0 FreeSans 224 0 0 0 N1END[0]
port 105 nsew signal input
flabel metal2 s 5814 0 5870 56 0 FreeSans 224 0 0 0 N1END[1]
port 106 nsew signal input
flabel metal2 s 5998 0 6054 56 0 FreeSans 224 0 0 0 N1END[2]
port 107 nsew signal input
flabel metal2 s 6182 0 6238 56 0 FreeSans 224 0 0 0 N1END[3]
port 108 nsew signal input
flabel metal2 s 7838 0 7894 56 0 FreeSans 224 0 0 0 N2END[0]
port 109 nsew signal input
flabel metal2 s 8022 0 8078 56 0 FreeSans 224 0 0 0 N2END[1]
port 110 nsew signal input
flabel metal2 s 8206 0 8262 56 0 FreeSans 224 0 0 0 N2END[2]
port 111 nsew signal input
flabel metal2 s 8390 0 8446 56 0 FreeSans 224 0 0 0 N2END[3]
port 112 nsew signal input
flabel metal2 s 8574 0 8630 56 0 FreeSans 224 0 0 0 N2END[4]
port 113 nsew signal input
flabel metal2 s 8758 0 8814 56 0 FreeSans 224 0 0 0 N2END[5]
port 114 nsew signal input
flabel metal2 s 8942 0 8998 56 0 FreeSans 224 0 0 0 N2END[6]
port 115 nsew signal input
flabel metal2 s 9126 0 9182 56 0 FreeSans 224 0 0 0 N2END[7]
port 116 nsew signal input
flabel metal2 s 6366 0 6422 56 0 FreeSans 224 0 0 0 N2MID[0]
port 117 nsew signal input
flabel metal2 s 6550 0 6606 56 0 FreeSans 224 0 0 0 N2MID[1]
port 118 nsew signal input
flabel metal2 s 6734 0 6790 56 0 FreeSans 224 0 0 0 N2MID[2]
port 119 nsew signal input
flabel metal2 s 6918 0 6974 56 0 FreeSans 224 0 0 0 N2MID[3]
port 120 nsew signal input
flabel metal2 s 7102 0 7158 56 0 FreeSans 224 0 0 0 N2MID[4]
port 121 nsew signal input
flabel metal2 s 7286 0 7342 56 0 FreeSans 224 0 0 0 N2MID[5]
port 122 nsew signal input
flabel metal2 s 7470 0 7526 56 0 FreeSans 224 0 0 0 N2MID[6]
port 123 nsew signal input
flabel metal2 s 7654 0 7710 56 0 FreeSans 224 0 0 0 N2MID[7]
port 124 nsew signal input
flabel metal2 s 9310 0 9366 56 0 FreeSans 224 0 0 0 N4END[0]
port 125 nsew signal input
flabel metal2 s 11150 0 11206 56 0 FreeSans 224 0 0 0 N4END[10]
port 126 nsew signal input
flabel metal2 s 11334 0 11390 56 0 FreeSans 224 0 0 0 N4END[11]
port 127 nsew signal input
flabel metal2 s 11518 0 11574 56 0 FreeSans 224 0 0 0 N4END[12]
port 128 nsew signal input
flabel metal2 s 11702 0 11758 56 0 FreeSans 224 0 0 0 N4END[13]
port 129 nsew signal input
flabel metal2 s 11886 0 11942 56 0 FreeSans 224 0 0 0 N4END[14]
port 130 nsew signal input
flabel metal2 s 12070 0 12126 56 0 FreeSans 224 0 0 0 N4END[15]
port 131 nsew signal input
flabel metal2 s 9494 0 9550 56 0 FreeSans 224 0 0 0 N4END[1]
port 132 nsew signal input
flabel metal2 s 9678 0 9734 56 0 FreeSans 224 0 0 0 N4END[2]
port 133 nsew signal input
flabel metal2 s 9862 0 9918 56 0 FreeSans 224 0 0 0 N4END[3]
port 134 nsew signal input
flabel metal2 s 10046 0 10102 56 0 FreeSans 224 0 0 0 N4END[4]
port 135 nsew signal input
flabel metal2 s 10230 0 10286 56 0 FreeSans 224 0 0 0 N4END[5]
port 136 nsew signal input
flabel metal2 s 10414 0 10470 56 0 FreeSans 224 0 0 0 N4END[6]
port 137 nsew signal input
flabel metal2 s 10598 0 10654 56 0 FreeSans 224 0 0 0 N4END[7]
port 138 nsew signal input
flabel metal2 s 10782 0 10838 56 0 FreeSans 224 0 0 0 N4END[8]
port 139 nsew signal input
flabel metal2 s 10966 0 11022 56 0 FreeSans 224 0 0 0 N4END[9]
port 140 nsew signal input
flabel metal2 s 12254 0 12310 56 0 FreeSans 224 0 0 0 NN4END[0]
port 141 nsew signal input
flabel metal2 s 14094 0 14150 56 0 FreeSans 224 0 0 0 NN4END[10]
port 142 nsew signal input
flabel metal2 s 14278 0 14334 56 0 FreeSans 224 0 0 0 NN4END[11]
port 143 nsew signal input
flabel metal2 s 14462 0 14518 56 0 FreeSans 224 0 0 0 NN4END[12]
port 144 nsew signal input
flabel metal2 s 14646 0 14702 56 0 FreeSans 224 0 0 0 NN4END[13]
port 145 nsew signal input
flabel metal2 s 14830 0 14886 56 0 FreeSans 224 0 0 0 NN4END[14]
port 146 nsew signal input
flabel metal2 s 15014 0 15070 56 0 FreeSans 224 0 0 0 NN4END[15]
port 147 nsew signal input
flabel metal2 s 12438 0 12494 56 0 FreeSans 224 0 0 0 NN4END[1]
port 148 nsew signal input
flabel metal2 s 12622 0 12678 56 0 FreeSans 224 0 0 0 NN4END[2]
port 149 nsew signal input
flabel metal2 s 12806 0 12862 56 0 FreeSans 224 0 0 0 NN4END[3]
port 150 nsew signal input
flabel metal2 s 12990 0 13046 56 0 FreeSans 224 0 0 0 NN4END[4]
port 151 nsew signal input
flabel metal2 s 13174 0 13230 56 0 FreeSans 224 0 0 0 NN4END[5]
port 152 nsew signal input
flabel metal2 s 13358 0 13414 56 0 FreeSans 224 0 0 0 NN4END[6]
port 153 nsew signal input
flabel metal2 s 13542 0 13598 56 0 FreeSans 224 0 0 0 NN4END[7]
port 154 nsew signal input
flabel metal2 s 13726 0 13782 56 0 FreeSans 224 0 0 0 NN4END[8]
port 155 nsew signal input
flabel metal2 s 13910 0 13966 56 0 FreeSans 224 0 0 0 NN4END[9]
port 156 nsew signal input
flabel metal2 s 15382 0 15438 56 0 FreeSans 224 0 0 0 S1BEG[0]
port 157 nsew signal output
flabel metal2 s 15566 0 15622 56 0 FreeSans 224 0 0 0 S1BEG[1]
port 158 nsew signal output
flabel metal2 s 15750 0 15806 56 0 FreeSans 224 0 0 0 S1BEG[2]
port 159 nsew signal output
flabel metal2 s 15934 0 15990 56 0 FreeSans 224 0 0 0 S1BEG[3]
port 160 nsew signal output
flabel metal2 s 16118 0 16174 56 0 FreeSans 224 0 0 0 S2BEG[0]
port 161 nsew signal output
flabel metal2 s 16302 0 16358 56 0 FreeSans 224 0 0 0 S2BEG[1]
port 162 nsew signal output
flabel metal2 s 16486 0 16542 56 0 FreeSans 224 0 0 0 S2BEG[2]
port 163 nsew signal output
flabel metal2 s 16670 0 16726 56 0 FreeSans 224 0 0 0 S2BEG[3]
port 164 nsew signal output
flabel metal2 s 16854 0 16910 56 0 FreeSans 224 0 0 0 S2BEG[4]
port 165 nsew signal output
flabel metal2 s 17038 0 17094 56 0 FreeSans 224 0 0 0 S2BEG[5]
port 166 nsew signal output
flabel metal2 s 17222 0 17278 56 0 FreeSans 224 0 0 0 S2BEG[6]
port 167 nsew signal output
flabel metal2 s 17406 0 17462 56 0 FreeSans 224 0 0 0 S2BEG[7]
port 168 nsew signal output
flabel metal2 s 17590 0 17646 56 0 FreeSans 224 0 0 0 S2BEGb[0]
port 169 nsew signal output
flabel metal2 s 17774 0 17830 56 0 FreeSans 224 0 0 0 S2BEGb[1]
port 170 nsew signal output
flabel metal2 s 17958 0 18014 56 0 FreeSans 224 0 0 0 S2BEGb[2]
port 171 nsew signal output
flabel metal2 s 18142 0 18198 56 0 FreeSans 224 0 0 0 S2BEGb[3]
port 172 nsew signal output
flabel metal2 s 18326 0 18382 56 0 FreeSans 224 0 0 0 S2BEGb[4]
port 173 nsew signal output
flabel metal2 s 18510 0 18566 56 0 FreeSans 224 0 0 0 S2BEGb[5]
port 174 nsew signal output
flabel metal2 s 18694 0 18750 56 0 FreeSans 224 0 0 0 S2BEGb[6]
port 175 nsew signal output
flabel metal2 s 18878 0 18934 56 0 FreeSans 224 0 0 0 S2BEGb[7]
port 176 nsew signal output
flabel metal2 s 19062 0 19118 56 0 FreeSans 224 0 0 0 S4BEG[0]
port 177 nsew signal output
flabel metal2 s 20902 0 20958 56 0 FreeSans 224 0 0 0 S4BEG[10]
port 178 nsew signal output
flabel metal2 s 21086 0 21142 56 0 FreeSans 224 0 0 0 S4BEG[11]
port 179 nsew signal output
flabel metal2 s 21270 0 21326 56 0 FreeSans 224 0 0 0 S4BEG[12]
port 180 nsew signal output
flabel metal2 s 21454 0 21510 56 0 FreeSans 224 0 0 0 S4BEG[13]
port 181 nsew signal output
flabel metal2 s 21638 0 21694 56 0 FreeSans 224 0 0 0 S4BEG[14]
port 182 nsew signal output
flabel metal2 s 21822 0 21878 56 0 FreeSans 224 0 0 0 S4BEG[15]
port 183 nsew signal output
flabel metal2 s 19246 0 19302 56 0 FreeSans 224 0 0 0 S4BEG[1]
port 184 nsew signal output
flabel metal2 s 19430 0 19486 56 0 FreeSans 224 0 0 0 S4BEG[2]
port 185 nsew signal output
flabel metal2 s 19614 0 19670 56 0 FreeSans 224 0 0 0 S4BEG[3]
port 186 nsew signal output
flabel metal2 s 19798 0 19854 56 0 FreeSans 224 0 0 0 S4BEG[4]
port 187 nsew signal output
flabel metal2 s 19982 0 20038 56 0 FreeSans 224 0 0 0 S4BEG[5]
port 188 nsew signal output
flabel metal2 s 20166 0 20222 56 0 FreeSans 224 0 0 0 S4BEG[6]
port 189 nsew signal output
flabel metal2 s 20350 0 20406 56 0 FreeSans 224 0 0 0 S4BEG[7]
port 190 nsew signal output
flabel metal2 s 20534 0 20590 56 0 FreeSans 224 0 0 0 S4BEG[8]
port 191 nsew signal output
flabel metal2 s 20718 0 20774 56 0 FreeSans 224 0 0 0 S4BEG[9]
port 192 nsew signal output
flabel metal2 s 22006 0 22062 56 0 FreeSans 224 0 0 0 SS4BEG[0]
port 193 nsew signal output
flabel metal2 s 23846 0 23902 56 0 FreeSans 224 0 0 0 SS4BEG[10]
port 194 nsew signal output
flabel metal2 s 24030 0 24086 56 0 FreeSans 224 0 0 0 SS4BEG[11]
port 195 nsew signal output
flabel metal2 s 24214 0 24270 56 0 FreeSans 224 0 0 0 SS4BEG[12]
port 196 nsew signal output
flabel metal2 s 24398 0 24454 56 0 FreeSans 224 0 0 0 SS4BEG[13]
port 197 nsew signal output
flabel metal2 s 24582 0 24638 56 0 FreeSans 224 0 0 0 SS4BEG[14]
port 198 nsew signal output
flabel metal2 s 24766 0 24822 56 0 FreeSans 224 0 0 0 SS4BEG[15]
port 199 nsew signal output
flabel metal2 s 22190 0 22246 56 0 FreeSans 224 0 0 0 SS4BEG[1]
port 200 nsew signal output
flabel metal2 s 22374 0 22430 56 0 FreeSans 224 0 0 0 SS4BEG[2]
port 201 nsew signal output
flabel metal2 s 22558 0 22614 56 0 FreeSans 224 0 0 0 SS4BEG[3]
port 202 nsew signal output
flabel metal2 s 22742 0 22798 56 0 FreeSans 224 0 0 0 SS4BEG[4]
port 203 nsew signal output
flabel metal2 s 22926 0 22982 56 0 FreeSans 224 0 0 0 SS4BEG[5]
port 204 nsew signal output
flabel metal2 s 23110 0 23166 56 0 FreeSans 224 0 0 0 SS4BEG[6]
port 205 nsew signal output
flabel metal2 s 23294 0 23350 56 0 FreeSans 224 0 0 0 SS4BEG[7]
port 206 nsew signal output
flabel metal2 s 23478 0 23534 56 0 FreeSans 224 0 0 0 SS4BEG[8]
port 207 nsew signal output
flabel metal2 s 23662 0 23718 56 0 FreeSans 224 0 0 0 SS4BEG[9]
port 208 nsew signal output
flabel metal2 s 24950 0 25006 56 0 FreeSans 224 0 0 0 UserCLK
port 209 nsew signal input
flabel metal2 s 1490 11096 1546 11152 0 FreeSans 224 0 0 0 UserCLKo
port 210 nsew signal output
flabel metal4 s 3004 0 3324 11152 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 3004 11092 3324 11152 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 9004 0 9324 11152 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 9004 0 9324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 9004 11092 9324 11152 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 15004 0 15324 11152 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 15004 0 15324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 15004 11092 15324 11152 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 21004 0 21324 11152 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 21004 0 21324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 21004 11092 21324 11152 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 27004 0 27324 11152 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 27004 0 27324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 27004 11092 27324 11152 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 33004 0 33324 11152 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 33004 0 33324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 33004 11092 33324 11152 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 1944 0 2264 11152 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 1944 11092 2264 11152 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 7944 0 8264 11152 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 7944 11092 8264 11152 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 13944 0 14264 11152 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 13944 0 14264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 13944 11092 14264 11152 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 19944 0 20264 11152 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 19944 0 20264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 19944 11092 20264 11152 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 25944 0 26264 11152 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 25944 0 26264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 25944 11092 26264 11152 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 31944 0 32264 11152 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 31944 0 32264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 31944 11092 32264 11152 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
rlabel metal1 17214 8704 17214 8704 0 VGND
rlabel metal1 17204 8160 17204 8160 0 VPWR
rlabel metal3 8900 1156 8900 1156 0 FrameData[0]
rlabel metal3 896 3876 896 3876 0 FrameData[10]
rlabel metal3 620 4148 620 4148 0 FrameData[11]
rlabel metal3 666 4420 666 4420 0 FrameData[12]
rlabel metal3 482 4692 482 4692 0 FrameData[13]
rlabel metal3 712 4964 712 4964 0 FrameData[14]
rlabel metal3 1402 5236 1402 5236 0 FrameData[15]
rlabel metal3 1448 5508 1448 5508 0 FrameData[16]
rlabel metal2 22310 6477 22310 6477 0 FrameData[17]
rlabel metal3 942 6052 942 6052 0 FrameData[18]
rlabel metal1 16836 6358 16836 6358 0 FrameData[19]
rlabel metal2 19458 1904 19458 1904 0 FrameData[1]
rlabel metal3 1494 6596 1494 6596 0 FrameData[20]
rlabel metal2 15778 5729 15778 5729 0 FrameData[21]
rlabel metal3 919 7140 919 7140 0 FrameData[22]
rlabel metal2 15410 5015 15410 5015 0 FrameData[23]
rlabel metal3 1494 7684 1494 7684 0 FrameData[24]
rlabel metal3 1356 7956 1356 7956 0 FrameData[25]
rlabel metal3 942 8228 942 8228 0 FrameData[26]
rlabel metal2 17066 7191 17066 7191 0 FrameData[27]
rlabel metal3 1448 8772 1448 8772 0 FrameData[28]
rlabel metal1 15042 5202 15042 5202 0 FrameData[29]
rlabel metal3 8440 1700 8440 1700 0 FrameData[2]
rlabel metal1 17020 5202 17020 5202 0 FrameData[30]
rlabel metal3 712 9588 712 9588 0 FrameData[31]
rlabel metal3 11016 1972 11016 1972 0 FrameData[3]
rlabel metal3 1494 2244 1494 2244 0 FrameData[4]
rlabel metal3 11752 2516 11752 2516 0 FrameData[5]
rlabel metal3 712 2788 712 2788 0 FrameData[6]
rlabel metal2 23598 3213 23598 3213 0 FrameData[7]
rlabel metal3 1494 3332 1494 3332 0 FrameData[8]
rlabel via2 20746 3587 20746 3587 0 FrameData[9]
rlabel metal3 33098 1156 33098 1156 0 FrameData_O[0]
rlabel metal3 33420 3876 33420 3876 0 FrameData_O[10]
rlabel metal3 33604 4148 33604 4148 0 FrameData_O[11]
rlabel metal3 33880 4420 33880 4420 0 FrameData_O[12]
rlabel metal3 33604 4692 33604 4692 0 FrameData_O[13]
rlabel metal3 33420 4964 33420 4964 0 FrameData_O[14]
rlabel metal3 33604 5236 33604 5236 0 FrameData_O[15]
rlabel metal3 33880 5508 33880 5508 0 FrameData_O[16]
rlabel metal3 33604 5780 33604 5780 0 FrameData_O[17]
rlabel metal3 33420 6052 33420 6052 0 FrameData_O[18]
rlabel metal3 33604 6324 33604 6324 0 FrameData_O[19]
rlabel metal2 31510 1853 31510 1853 0 FrameData_O[1]
rlabel metal1 32522 6664 32522 6664 0 FrameData_O[20]
rlabel metal2 32890 6749 32890 6749 0 FrameData_O[21]
rlabel metal3 33604 7140 33604 7140 0 FrameData_O[22]
rlabel metal3 33420 7412 33420 7412 0 FrameData_O[23]
rlabel metal3 33972 7684 33972 7684 0 FrameData_O[24]
rlabel metal3 33420 7956 33420 7956 0 FrameData_O[25]
rlabel metal3 33696 8228 33696 8228 0 FrameData_O[26]
rlabel metal1 32246 8058 32246 8058 0 FrameData_O[27]
rlabel metal1 32982 7514 32982 7514 0 FrameData_O[28]
rlabel metal2 31786 8551 31786 8551 0 FrameData_O[29]
rlabel metal3 33374 1700 33374 1700 0 FrameData_O[2]
rlabel metal2 31142 8959 31142 8959 0 FrameData_O[30]
rlabel metal2 31418 8823 31418 8823 0 FrameData_O[31]
rlabel metal2 31142 2125 31142 2125 0 FrameData_O[3]
rlabel metal3 33880 2244 33880 2244 0 FrameData_O[4]
rlabel metal3 33604 2516 33604 2516 0 FrameData_O[5]
rlabel metal3 33420 2788 33420 2788 0 FrameData_O[6]
rlabel metal3 33604 3060 33604 3060 0 FrameData_O[7]
rlabel metal3 33880 3332 33880 3332 0 FrameData_O[8]
rlabel metal3 33604 3604 33604 3604 0 FrameData_O[9]
rlabel metal1 9568 7378 9568 7378 0 FrameStrobe[0]
rlabel metal2 27002 667 27002 667 0 FrameStrobe[10]
rlabel metal2 27186 718 27186 718 0 FrameStrobe[11]
rlabel metal2 27370 820 27370 820 0 FrameStrobe[12]
rlabel metal2 27554 735 27554 735 0 FrameStrobe[13]
rlabel metal2 27738 922 27738 922 0 FrameStrobe[14]
rlabel metal2 27922 55 27922 55 0 FrameStrobe[15]
rlabel metal1 28520 6766 28520 6766 0 FrameStrobe[16]
rlabel metal2 28290 718 28290 718 0 FrameStrobe[17]
rlabel metal2 28474 786 28474 786 0 FrameStrobe[18]
rlabel metal1 28704 5202 28704 5202 0 FrameStrobe[19]
rlabel metal2 12374 7548 12374 7548 0 FrameStrobe[1]
rlabel metal1 14858 7378 14858 7378 0 FrameStrobe[2]
rlabel metal2 14398 7616 14398 7616 0 FrameStrobe[3]
rlabel metal2 25898 395 25898 395 0 FrameStrobe[4]
rlabel metal2 26082 1279 26082 1279 0 FrameStrobe[5]
rlabel metal2 26266 55 26266 55 0 FrameStrobe[6]
rlabel metal1 26358 6766 26358 6766 0 FrameStrobe[7]
rlabel via2 26634 55 26634 55 0 FrameStrobe[8]
rlabel metal2 26818 718 26818 718 0 FrameStrobe[9]
rlabel metal1 3082 8602 3082 8602 0 FrameStrobe_O[0]
rlabel metal1 18814 8602 18814 8602 0 FrameStrobe_O[10]
rlabel metal1 20378 8602 20378 8602 0 FrameStrobe_O[11]
rlabel metal1 21942 8602 21942 8602 0 FrameStrobe_O[12]
rlabel metal1 23506 8602 23506 8602 0 FrameStrobe_O[13]
rlabel metal1 25116 8602 25116 8602 0 FrameStrobe_O[14]
rlabel metal1 26818 8602 26818 8602 0 FrameStrobe_O[15]
rlabel metal1 28198 8602 28198 8602 0 FrameStrobe_O[16]
rlabel metal1 29808 8602 29808 8602 0 FrameStrobe_O[17]
rlabel metal1 31372 8602 31372 8602 0 FrameStrobe_O[18]
rlabel metal1 32844 8602 32844 8602 0 FrameStrobe_O[19]
rlabel metal1 4738 8602 4738 8602 0 FrameStrobe_O[1]
rlabel metal1 6348 8602 6348 8602 0 FrameStrobe_O[2]
rlabel metal1 7866 8602 7866 8602 0 FrameStrobe_O[3]
rlabel metal1 9476 8602 9476 8602 0 FrameStrobe_O[4]
rlabel metal1 10994 8330 10994 8330 0 FrameStrobe_O[5]
rlabel metal1 12558 8602 12558 8602 0 FrameStrobe_O[6]
rlabel metal1 14122 8602 14122 8602 0 FrameStrobe_O[7]
rlabel metal1 15686 8602 15686 8602 0 FrameStrobe_O[8]
rlabel metal1 17250 8602 17250 8602 0 FrameStrobe_O[9]
rlabel metal2 5658 1976 5658 1976 0 N1END[0]
rlabel metal2 5842 2316 5842 2316 0 N1END[1]
rlabel metal2 6026 2282 6026 2282 0 N1END[2]
rlabel metal2 6210 2350 6210 2350 0 N1END[3]
rlabel metal2 7866 123 7866 123 0 N2END[0]
rlabel metal2 8050 1007 8050 1007 0 N2END[1]
rlabel metal2 8234 1075 8234 1075 0 N2END[2]
rlabel metal2 8418 1806 8418 1806 0 N2END[3]
rlabel metal2 8602 2078 8602 2078 0 N2END[4]
rlabel metal2 8786 1772 8786 1772 0 N2END[5]
rlabel metal2 8970 55 8970 55 0 N2END[6]
rlabel metal2 6578 3774 6578 3774 0 N2END[7]
rlabel metal2 6394 2078 6394 2078 0 N2MID[0]
rlabel metal2 6578 55 6578 55 0 N2MID[1]
rlabel metal2 6762 1874 6762 1874 0 N2MID[2]
rlabel metal2 3450 3876 3450 3876 0 N2MID[3]
rlabel metal2 7130 1772 7130 1772 0 N2MID[4]
rlabel metal2 2898 3808 2898 3808 0 N2MID[5]
rlabel metal2 4554 2227 4554 2227 0 N2MID[6]
rlabel metal2 4922 1751 4922 1751 0 N2MID[7]
rlabel metal2 9338 684 9338 684 0 N4END[0]
rlabel metal2 11178 2282 11178 2282 0 N4END[10]
rlabel metal2 11362 2316 11362 2316 0 N4END[11]
rlabel metal2 11546 2350 11546 2350 0 N4END[12]
rlabel metal2 11730 2384 11730 2384 0 N4END[13]
rlabel metal2 11914 55 11914 55 0 N4END[14]
rlabel metal2 12098 2282 12098 2282 0 N4END[15]
rlabel metal2 9522 650 9522 650 0 N4END[1]
rlabel metal2 9706 2010 9706 2010 0 N4END[2]
rlabel metal2 9890 1075 9890 1075 0 N4END[3]
rlabel metal2 10074 2622 10074 2622 0 N4END[4]
rlabel metal2 10258 1160 10258 1160 0 N4END[5]
rlabel metal2 10442 1228 10442 1228 0 N4END[6]
rlabel metal2 10626 1432 10626 1432 0 N4END[7]
rlabel metal2 10810 2146 10810 2146 0 N4END[8]
rlabel metal2 10994 2418 10994 2418 0 N4END[9]
rlabel metal2 12282 208 12282 208 0 NN4END[0]
rlabel metal2 14122 55 14122 55 0 NN4END[10]
rlabel metal2 14306 55 14306 55 0 NN4END[11]
rlabel metal2 14490 820 14490 820 0 NN4END[12]
rlabel metal2 14674 55 14674 55 0 NN4END[13]
rlabel metal2 14858 276 14858 276 0 NN4END[14]
rlabel metal2 15042 140 15042 140 0 NN4END[15]
rlabel metal2 12466 1211 12466 1211 0 NN4END[1]
rlabel metal2 12650 140 12650 140 0 NN4END[2]
rlabel metal2 12834 106 12834 106 0 NN4END[3]
rlabel metal2 13018 123 13018 123 0 NN4END[4]
rlabel metal2 13202 174 13202 174 0 NN4END[5]
rlabel metal2 13386 191 13386 191 0 NN4END[6]
rlabel metal2 13570 259 13570 259 0 NN4END[7]
rlabel metal2 13754 327 13754 327 0 NN4END[8]
rlabel metal2 13938 123 13938 123 0 NN4END[9]
rlabel metal1 15548 2822 15548 2822 0 S1BEG[0]
rlabel metal2 15594 1296 15594 1296 0 S1BEG[1]
rlabel metal1 15916 2822 15916 2822 0 S1BEG[2]
rlabel metal2 15962 1194 15962 1194 0 S1BEG[3]
rlabel metal1 16284 2822 16284 2822 0 S2BEG[0]
rlabel metal2 16330 1160 16330 1160 0 S2BEG[1]
rlabel metal2 16514 1296 16514 1296 0 S2BEG[2]
rlabel metal1 16836 2822 16836 2822 0 S2BEG[3]
rlabel metal2 16882 1160 16882 1160 0 S2BEG[4]
rlabel metal1 17204 2822 17204 2822 0 S2BEG[5]
rlabel metal2 17250 1160 17250 1160 0 S2BEG[6]
rlabel metal1 17572 2822 17572 2822 0 S2BEG[7]
rlabel metal2 17618 1160 17618 1160 0 S2BEGb[0]
rlabel metal2 17802 1160 17802 1160 0 S2BEGb[1]
rlabel metal2 17986 1160 17986 1160 0 S2BEGb[2]
rlabel metal2 18170 1296 18170 1296 0 S2BEGb[3]
rlabel metal2 18354 1160 18354 1160 0 S2BEGb[4]
rlabel metal2 18538 1330 18538 1330 0 S2BEGb[5]
rlabel metal2 18722 1160 18722 1160 0 S2BEGb[6]
rlabel metal1 19044 2822 19044 2822 0 S2BEGb[7]
rlabel metal2 19090 1194 19090 1194 0 S4BEG[0]
rlabel metal2 20930 1296 20930 1296 0 S4BEG[10]
rlabel metal2 21114 718 21114 718 0 S4BEG[11]
rlabel metal2 21298 55 21298 55 0 S4BEG[12]
rlabel metal2 21482 1194 21482 1194 0 S4BEG[13]
rlabel metal2 21666 1466 21666 1466 0 S4BEG[14]
rlabel metal2 21850 1330 21850 1330 0 S4BEG[15]
rlabel metal1 19412 2822 19412 2822 0 S4BEG[1]
rlabel metal2 19458 55 19458 55 0 S4BEG[2]
rlabel metal1 19780 2822 19780 2822 0 S4BEG[3]
rlabel metal2 19826 55 19826 55 0 S4BEG[4]
rlabel metal2 20010 55 20010 55 0 S4BEG[5]
rlabel metal2 20194 1330 20194 1330 0 S4BEG[6]
rlabel metal1 20516 2822 20516 2822 0 S4BEG[7]
rlabel metal1 20792 2890 20792 2890 0 S4BEG[8]
rlabel metal1 21068 2822 21068 2822 0 S4BEG[9]
rlabel metal2 22034 1602 22034 1602 0 SS4BEG[0]
rlabel metal2 23874 1194 23874 1194 0 SS4BEG[10]
rlabel metal1 24472 2890 24472 2890 0 SS4BEG[11]
rlabel metal2 24242 1330 24242 1330 0 SS4BEG[12]
rlabel metal1 24702 2822 24702 2822 0 SS4BEG[13]
rlabel metal2 24610 1160 24610 1160 0 SS4BEG[14]
rlabel metal1 25208 3162 25208 3162 0 SS4BEG[15]
rlabel metal2 22218 1296 22218 1296 0 SS4BEG[1]
rlabel metal2 22402 55 22402 55 0 SS4BEG[2]
rlabel metal2 22586 55 22586 55 0 SS4BEG[3]
rlabel metal1 23092 2822 23092 2822 0 SS4BEG[4]
rlabel metal1 23368 2958 23368 2958 0 SS4BEG[5]
rlabel metal2 23138 55 23138 55 0 SS4BEG[6]
rlabel metal1 23414 2890 23414 2890 0 SS4BEG[7]
rlabel metal2 23506 1296 23506 1296 0 SS4BEG[8]
rlabel metal1 24104 3162 24104 3162 0 SS4BEG[9]
rlabel metal1 11270 7344 11270 7344 0 UserCLK
rlabel metal1 1564 8602 1564 8602 0 UserCLKo
rlabel metal1 18676 3366 18676 3366 0 net1
rlabel metal2 32338 5814 32338 5814 0 net10
rlabel metal2 23966 3536 23966 3536 0 net100
rlabel metal1 24610 2414 24610 2414 0 net101
rlabel metal1 24334 3060 24334 3060 0 net102
rlabel metal1 25208 2414 25208 2414 0 net103
rlabel metal2 24702 3502 24702 3502 0 net104
rlabel metal1 1794 8500 1794 8500 0 net105
rlabel metal1 32706 6222 32706 6222 0 net11
rlabel metal1 21206 3604 21206 3604 0 net12
rlabel metal2 31786 5712 31786 5712 0 net13
rlabel metal1 32430 6698 32430 6698 0 net14
rlabel metal1 32706 7344 32706 7344 0 net15
rlabel metal1 32338 7922 32338 7922 0 net16
rlabel metal1 32706 7820 32706 7820 0 net17
rlabel metal1 32338 8432 32338 8432 0 net18
rlabel metal2 20470 6256 20470 6256 0 net19
rlabel metal2 30590 5644 30590 5644 0 net2
rlabel metal1 17618 5610 17618 5610 0 net20
rlabel metal1 19918 5576 19918 5576 0 net21
rlabel metal2 15594 5882 15594 5882 0 net22
rlabel metal1 21758 3400 21758 3400 0 net23
rlabel metal1 17296 5066 17296 5066 0 net24
rlabel metal1 21390 6664 21390 6664 0 net25
rlabel metal1 26542 1938 26542 1938 0 net26
rlabel metal2 32338 1938 32338 1938 0 net27
rlabel metal1 32706 2516 32706 2516 0 net28
rlabel metal1 32338 3060 32338 3060 0 net29
rlabel metal1 32706 4080 32706 4080 0 net3
rlabel metal1 32706 2958 32706 2958 0 net30
rlabel metal1 32338 3468 32338 3468 0 net31
rlabel metal1 32706 3536 32706 3536 0 net32
rlabel metal2 5566 7888 5566 7888 0 net33
rlabel metal1 19090 8500 19090 8500 0 net34
rlabel metal2 20654 8636 20654 8636 0 net35
rlabel metal2 29486 7922 29486 7922 0 net36
rlabel metal1 30912 7514 30912 7514 0 net37
rlabel metal2 24886 7548 24886 7548 0 net38
rlabel metal2 28014 7990 28014 7990 0 net39
rlabel metal1 32108 4590 32108 4590 0 net4
rlabel metal2 28750 7548 28750 7548 0 net40
rlabel metal2 29762 7446 29762 7446 0 net41
rlabel metal1 31188 5882 31188 5882 0 net42
rlabel metal1 32568 8466 32568 8466 0 net43
rlabel metal1 5014 8398 5014 8398 0 net44
rlabel metal2 8050 8636 8050 8636 0 net45
rlabel metal1 11178 8296 11178 8296 0 net46
rlabel metal2 24794 7888 24794 7888 0 net47
rlabel metal2 28290 8194 28290 8194 0 net48
rlabel metal2 12834 8738 12834 8738 0 net49
rlabel metal1 32706 4692 32706 4692 0 net5
rlabel metal2 14398 8772 14398 8772 0 net50
rlabel metal2 19458 7344 19458 7344 0 net51
rlabel metal2 19734 7514 19734 7514 0 net52
rlabel metal2 3174 4998 3174 4998 0 net53
rlabel metal2 3450 5032 3450 5032 0 net54
rlabel metal2 10166 3808 10166 3808 0 net55
rlabel metal2 4186 3196 4186 3196 0 net56
rlabel metal2 2714 3570 2714 3570 0 net57
rlabel metal2 2806 3264 2806 3264 0 net58
rlabel metal2 3542 3196 3542 3196 0 net59
rlabel metal1 32338 5168 32338 5168 0 net6
rlabel metal2 2530 3417 2530 3417 0 net60
rlabel metal2 3634 3264 3634 3264 0 net61
rlabel metal2 3910 3434 3910 3434 0 net62
rlabel metal2 4462 2788 4462 2788 0 net63
rlabel metal1 7406 4012 7406 4012 0 net64
rlabel metal2 7222 2890 7222 2890 0 net65
rlabel metal2 7406 5032 7406 5032 0 net66
rlabel metal2 7406 2550 7406 2550 0 net67
rlabel metal2 7038 3944 7038 3944 0 net68
rlabel metal2 7498 2958 7498 2958 0 net69
rlabel metal1 32706 5236 32706 5236 0 net7
rlabel metal2 13662 3706 13662 3706 0 net70
rlabel metal2 8326 2312 8326 2312 0 net71
rlabel metal2 7682 3808 7682 3808 0 net72
rlabel metal1 18216 2074 18216 2074 0 net73
rlabel metal1 21804 2414 21804 2414 0 net74
rlabel metal1 21620 2482 21620 2482 0 net75
rlabel metal2 21850 3536 21850 3536 0 net76
rlabel metal1 16652 1462 16652 1462 0 net77
rlabel metal2 22310 3502 22310 3502 0 net78
rlabel metal1 15502 3910 15502 3910 0 net79
rlabel metal2 24150 7208 24150 7208 0 net8
rlabel metal1 19320 3026 19320 3026 0 net80
rlabel metal1 19918 2482 19918 2482 0 net81
rlabel metal2 11270 4318 11270 4318 0 net82
rlabel metal2 11638 4573 11638 4573 0 net83
rlabel metal1 20102 3060 20102 3060 0 net84
rlabel metal2 12098 4896 12098 4896 0 net85
rlabel metal2 20470 3638 20470 3638 0 net86
rlabel metal2 17618 3264 17618 3264 0 net87
rlabel metal1 21206 2992 21206 2992 0 net88
rlabel metal2 22862 3570 22862 3570 0 net89
rlabel metal1 32706 5712 32706 5712 0 net9
rlabel metal2 27784 2652 27784 2652 0 net90
rlabel metal2 25070 3230 25070 3230 0 net91
rlabel metal1 26312 2482 26312 2482 0 net92
rlabel viali 25438 3028 25438 3028 0 net93
rlabel metal1 26450 2414 26450 2414 0 net94
rlabel metal2 25806 3196 25806 3196 0 net95
rlabel metal1 25898 2074 25898 2074 0 net96
rlabel metal2 23230 3876 23230 3876 0 net97
rlabel metal2 23966 2465 23966 2465 0 net98
rlabel metal1 23736 3026 23736 3026 0 net99
<< properties >>
string FIXED_BBOX 0 0 34408 11152
<< end >>
